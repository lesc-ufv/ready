module omega256x256_8_0_1 #
(
  parameter WIDTH = 16,
  parameter PIPE_EXTRA = 0
)
(
  input clk,
  input rst,
  input en,
  input [64-1:0] net_conf_bus_in,
  input [WIDTH-1:0] in0,
  input [WIDTH-1:0] in1,
  input [WIDTH-1:0] in2,
  input [WIDTH-1:0] in3,
  input [WIDTH-1:0] in4,
  input [WIDTH-1:0] in5,
  input [WIDTH-1:0] in6,
  input [WIDTH-1:0] in7,
  input [WIDTH-1:0] in8,
  input [WIDTH-1:0] in9,
  input [WIDTH-1:0] in10,
  input [WIDTH-1:0] in11,
  input [WIDTH-1:0] in12,
  input [WIDTH-1:0] in13,
  input [WIDTH-1:0] in14,
  input [WIDTH-1:0] in15,
  input [WIDTH-1:0] in16,
  input [WIDTH-1:0] in17,
  input [WIDTH-1:0] in18,
  input [WIDTH-1:0] in19,
  input [WIDTH-1:0] in20,
  input [WIDTH-1:0] in21,
  input [WIDTH-1:0] in22,
  input [WIDTH-1:0] in23,
  input [WIDTH-1:0] in24,
  input [WIDTH-1:0] in25,
  input [WIDTH-1:0] in26,
  input [WIDTH-1:0] in27,
  input [WIDTH-1:0] in28,
  input [WIDTH-1:0] in29,
  input [WIDTH-1:0] in30,
  input [WIDTH-1:0] in31,
  input [WIDTH-1:0] in32,
  input [WIDTH-1:0] in33,
  input [WIDTH-1:0] in34,
  input [WIDTH-1:0] in35,
  input [WIDTH-1:0] in36,
  input [WIDTH-1:0] in37,
  input [WIDTH-1:0] in38,
  input [WIDTH-1:0] in39,
  input [WIDTH-1:0] in40,
  input [WIDTH-1:0] in41,
  input [WIDTH-1:0] in42,
  input [WIDTH-1:0] in43,
  input [WIDTH-1:0] in44,
  input [WIDTH-1:0] in45,
  input [WIDTH-1:0] in46,
  input [WIDTH-1:0] in47,
  input [WIDTH-1:0] in48,
  input [WIDTH-1:0] in49,
  input [WIDTH-1:0] in50,
  input [WIDTH-1:0] in51,
  input [WIDTH-1:0] in52,
  input [WIDTH-1:0] in53,
  input [WIDTH-1:0] in54,
  input [WIDTH-1:0] in55,
  input [WIDTH-1:0] in56,
  input [WIDTH-1:0] in57,
  input [WIDTH-1:0] in58,
  input [WIDTH-1:0] in59,
  input [WIDTH-1:0] in60,
  input [WIDTH-1:0] in61,
  input [WIDTH-1:0] in62,
  input [WIDTH-1:0] in63,
  input [WIDTH-1:0] in64,
  input [WIDTH-1:0] in65,
  input [WIDTH-1:0] in66,
  input [WIDTH-1:0] in67,
  input [WIDTH-1:0] in68,
  input [WIDTH-1:0] in69,
  input [WIDTH-1:0] in70,
  input [WIDTH-1:0] in71,
  input [WIDTH-1:0] in72,
  input [WIDTH-1:0] in73,
  input [WIDTH-1:0] in74,
  input [WIDTH-1:0] in75,
  input [WIDTH-1:0] in76,
  input [WIDTH-1:0] in77,
  input [WIDTH-1:0] in78,
  input [WIDTH-1:0] in79,
  input [WIDTH-1:0] in80,
  input [WIDTH-1:0] in81,
  input [WIDTH-1:0] in82,
  input [WIDTH-1:0] in83,
  input [WIDTH-1:0] in84,
  input [WIDTH-1:0] in85,
  input [WIDTH-1:0] in86,
  input [WIDTH-1:0] in87,
  input [WIDTH-1:0] in88,
  input [WIDTH-1:0] in89,
  input [WIDTH-1:0] in90,
  input [WIDTH-1:0] in91,
  input [WIDTH-1:0] in92,
  input [WIDTH-1:0] in93,
  input [WIDTH-1:0] in94,
  input [WIDTH-1:0] in95,
  input [WIDTH-1:0] in96,
  input [WIDTH-1:0] in97,
  input [WIDTH-1:0] in98,
  input [WIDTH-1:0] in99,
  input [WIDTH-1:0] in100,
  input [WIDTH-1:0] in101,
  input [WIDTH-1:0] in102,
  input [WIDTH-1:0] in103,
  input [WIDTH-1:0] in104,
  input [WIDTH-1:0] in105,
  input [WIDTH-1:0] in106,
  input [WIDTH-1:0] in107,
  input [WIDTH-1:0] in108,
  input [WIDTH-1:0] in109,
  input [WIDTH-1:0] in110,
  input [WIDTH-1:0] in111,
  input [WIDTH-1:0] in112,
  input [WIDTH-1:0] in113,
  input [WIDTH-1:0] in114,
  input [WIDTH-1:0] in115,
  input [WIDTH-1:0] in116,
  input [WIDTH-1:0] in117,
  input [WIDTH-1:0] in118,
  input [WIDTH-1:0] in119,
  input [WIDTH-1:0] in120,
  input [WIDTH-1:0] in121,
  input [WIDTH-1:0] in122,
  input [WIDTH-1:0] in123,
  input [WIDTH-1:0] in124,
  input [WIDTH-1:0] in125,
  input [WIDTH-1:0] in126,
  input [WIDTH-1:0] in127,
  input [WIDTH-1:0] in128,
  input [WIDTH-1:0] in129,
  input [WIDTH-1:0] in130,
  input [WIDTH-1:0] in131,
  input [WIDTH-1:0] in132,
  input [WIDTH-1:0] in133,
  input [WIDTH-1:0] in134,
  input [WIDTH-1:0] in135,
  input [WIDTH-1:0] in136,
  input [WIDTH-1:0] in137,
  input [WIDTH-1:0] in138,
  input [WIDTH-1:0] in139,
  input [WIDTH-1:0] in140,
  input [WIDTH-1:0] in141,
  input [WIDTH-1:0] in142,
  input [WIDTH-1:0] in143,
  input [WIDTH-1:0] in144,
  input [WIDTH-1:0] in145,
  input [WIDTH-1:0] in146,
  input [WIDTH-1:0] in147,
  input [WIDTH-1:0] in148,
  input [WIDTH-1:0] in149,
  input [WIDTH-1:0] in150,
  input [WIDTH-1:0] in151,
  input [WIDTH-1:0] in152,
  input [WIDTH-1:0] in153,
  input [WIDTH-1:0] in154,
  input [WIDTH-1:0] in155,
  input [WIDTH-1:0] in156,
  input [WIDTH-1:0] in157,
  input [WIDTH-1:0] in158,
  input [WIDTH-1:0] in159,
  input [WIDTH-1:0] in160,
  input [WIDTH-1:0] in161,
  input [WIDTH-1:0] in162,
  input [WIDTH-1:0] in163,
  input [WIDTH-1:0] in164,
  input [WIDTH-1:0] in165,
  input [WIDTH-1:0] in166,
  input [WIDTH-1:0] in167,
  input [WIDTH-1:0] in168,
  input [WIDTH-1:0] in169,
  input [WIDTH-1:0] in170,
  input [WIDTH-1:0] in171,
  input [WIDTH-1:0] in172,
  input [WIDTH-1:0] in173,
  input [WIDTH-1:0] in174,
  input [WIDTH-1:0] in175,
  input [WIDTH-1:0] in176,
  input [WIDTH-1:0] in177,
  input [WIDTH-1:0] in178,
  input [WIDTH-1:0] in179,
  input [WIDTH-1:0] in180,
  input [WIDTH-1:0] in181,
  input [WIDTH-1:0] in182,
  input [WIDTH-1:0] in183,
  input [WIDTH-1:0] in184,
  input [WIDTH-1:0] in185,
  input [WIDTH-1:0] in186,
  input [WIDTH-1:0] in187,
  input [WIDTH-1:0] in188,
  input [WIDTH-1:0] in189,
  input [WIDTH-1:0] in190,
  input [WIDTH-1:0] in191,
  input [WIDTH-1:0] in192,
  input [WIDTH-1:0] in193,
  input [WIDTH-1:0] in194,
  input [WIDTH-1:0] in195,
  input [WIDTH-1:0] in196,
  input [WIDTH-1:0] in197,
  input [WIDTH-1:0] in198,
  input [WIDTH-1:0] in199,
  input [WIDTH-1:0] in200,
  input [WIDTH-1:0] in201,
  input [WIDTH-1:0] in202,
  input [WIDTH-1:0] in203,
  input [WIDTH-1:0] in204,
  input [WIDTH-1:0] in205,
  input [WIDTH-1:0] in206,
  input [WIDTH-1:0] in207,
  input [WIDTH-1:0] in208,
  input [WIDTH-1:0] in209,
  input [WIDTH-1:0] in210,
  input [WIDTH-1:0] in211,
  input [WIDTH-1:0] in212,
  input [WIDTH-1:0] in213,
  input [WIDTH-1:0] in214,
  input [WIDTH-1:0] in215,
  input [WIDTH-1:0] in216,
  input [WIDTH-1:0] in217,
  input [WIDTH-1:0] in218,
  input [WIDTH-1:0] in219,
  input [WIDTH-1:0] in220,
  input [WIDTH-1:0] in221,
  input [WIDTH-1:0] in222,
  input [WIDTH-1:0] in223,
  input [WIDTH-1:0] in224,
  input [WIDTH-1:0] in225,
  input [WIDTH-1:0] in226,
  input [WIDTH-1:0] in227,
  input [WIDTH-1:0] in228,
  input [WIDTH-1:0] in229,
  input [WIDTH-1:0] in230,
  input [WIDTH-1:0] in231,
  input [WIDTH-1:0] in232,
  input [WIDTH-1:0] in233,
  input [WIDTH-1:0] in234,
  input [WIDTH-1:0] in235,
  input [WIDTH-1:0] in236,
  input [WIDTH-1:0] in237,
  input [WIDTH-1:0] in238,
  input [WIDTH-1:0] in239,
  input [WIDTH-1:0] in240,
  input [WIDTH-1:0] in241,
  input [WIDTH-1:0] in242,
  input [WIDTH-1:0] in243,
  input [WIDTH-1:0] in244,
  input [WIDTH-1:0] in245,
  input [WIDTH-1:0] in246,
  input [WIDTH-1:0] in247,
  input [WIDTH-1:0] in248,
  input [WIDTH-1:0] in249,
  input [WIDTH-1:0] in250,
  input [WIDTH-1:0] in251,
  input [WIDTH-1:0] in252,
  input [WIDTH-1:0] in253,
  input [WIDTH-1:0] in254,
  input [WIDTH-1:0] in255,
  output [WIDTH-1:0] out0,
  output [WIDTH-1:0] out1,
  output [WIDTH-1:0] out2,
  output [WIDTH-1:0] out3,
  output [WIDTH-1:0] out4,
  output [WIDTH-1:0] out5,
  output [WIDTH-1:0] out6,
  output [WIDTH-1:0] out7,
  output [WIDTH-1:0] out8,
  output [WIDTH-1:0] out9,
  output [WIDTH-1:0] out10,
  output [WIDTH-1:0] out11,
  output [WIDTH-1:0] out12,
  output [WIDTH-1:0] out13,
  output [WIDTH-1:0] out14,
  output [WIDTH-1:0] out15,
  output [WIDTH-1:0] out16,
  output [WIDTH-1:0] out17,
  output [WIDTH-1:0] out18,
  output [WIDTH-1:0] out19,
  output [WIDTH-1:0] out20,
  output [WIDTH-1:0] out21,
  output [WIDTH-1:0] out22,
  output [WIDTH-1:0] out23,
  output [WIDTH-1:0] out24,
  output [WIDTH-1:0] out25,
  output [WIDTH-1:0] out26,
  output [WIDTH-1:0] out27,
  output [WIDTH-1:0] out28,
  output [WIDTH-1:0] out29,
  output [WIDTH-1:0] out30,
  output [WIDTH-1:0] out31,
  output [WIDTH-1:0] out32,
  output [WIDTH-1:0] out33,
  output [WIDTH-1:0] out34,
  output [WIDTH-1:0] out35,
  output [WIDTH-1:0] out36,
  output [WIDTH-1:0] out37,
  output [WIDTH-1:0] out38,
  output [WIDTH-1:0] out39,
  output [WIDTH-1:0] out40,
  output [WIDTH-1:0] out41,
  output [WIDTH-1:0] out42,
  output [WIDTH-1:0] out43,
  output [WIDTH-1:0] out44,
  output [WIDTH-1:0] out45,
  output [WIDTH-1:0] out46,
  output [WIDTH-1:0] out47,
  output [WIDTH-1:0] out48,
  output [WIDTH-1:0] out49,
  output [WIDTH-1:0] out50,
  output [WIDTH-1:0] out51,
  output [WIDTH-1:0] out52,
  output [WIDTH-1:0] out53,
  output [WIDTH-1:0] out54,
  output [WIDTH-1:0] out55,
  output [WIDTH-1:0] out56,
  output [WIDTH-1:0] out57,
  output [WIDTH-1:0] out58,
  output [WIDTH-1:0] out59,
  output [WIDTH-1:0] out60,
  output [WIDTH-1:0] out61,
  output [WIDTH-1:0] out62,
  output [WIDTH-1:0] out63,
  output [WIDTH-1:0] out64,
  output [WIDTH-1:0] out65,
  output [WIDTH-1:0] out66,
  output [WIDTH-1:0] out67,
  output [WIDTH-1:0] out68,
  output [WIDTH-1:0] out69,
  output [WIDTH-1:0] out70,
  output [WIDTH-1:0] out71,
  output [WIDTH-1:0] out72,
  output [WIDTH-1:0] out73,
  output [WIDTH-1:0] out74,
  output [WIDTH-1:0] out75,
  output [WIDTH-1:0] out76,
  output [WIDTH-1:0] out77,
  output [WIDTH-1:0] out78,
  output [WIDTH-1:0] out79,
  output [WIDTH-1:0] out80,
  output [WIDTH-1:0] out81,
  output [WIDTH-1:0] out82,
  output [WIDTH-1:0] out83,
  output [WIDTH-1:0] out84,
  output [WIDTH-1:0] out85,
  output [WIDTH-1:0] out86,
  output [WIDTH-1:0] out87,
  output [WIDTH-1:0] out88,
  output [WIDTH-1:0] out89,
  output [WIDTH-1:0] out90,
  output [WIDTH-1:0] out91,
  output [WIDTH-1:0] out92,
  output [WIDTH-1:0] out93,
  output [WIDTH-1:0] out94,
  output [WIDTH-1:0] out95,
  output [WIDTH-1:0] out96,
  output [WIDTH-1:0] out97,
  output [WIDTH-1:0] out98,
  output [WIDTH-1:0] out99,
  output [WIDTH-1:0] out100,
  output [WIDTH-1:0] out101,
  output [WIDTH-1:0] out102,
  output [WIDTH-1:0] out103,
  output [WIDTH-1:0] out104,
  output [WIDTH-1:0] out105,
  output [WIDTH-1:0] out106,
  output [WIDTH-1:0] out107,
  output [WIDTH-1:0] out108,
  output [WIDTH-1:0] out109,
  output [WIDTH-1:0] out110,
  output [WIDTH-1:0] out111,
  output [WIDTH-1:0] out112,
  output [WIDTH-1:0] out113,
  output [WIDTH-1:0] out114,
  output [WIDTH-1:0] out115,
  output [WIDTH-1:0] out116,
  output [WIDTH-1:0] out117,
  output [WIDTH-1:0] out118,
  output [WIDTH-1:0] out119,
  output [WIDTH-1:0] out120,
  output [WIDTH-1:0] out121,
  output [WIDTH-1:0] out122,
  output [WIDTH-1:0] out123,
  output [WIDTH-1:0] out124,
  output [WIDTH-1:0] out125,
  output [WIDTH-1:0] out126,
  output [WIDTH-1:0] out127,
  output [WIDTH-1:0] out128,
  output [WIDTH-1:0] out129,
  output [WIDTH-1:0] out130,
  output [WIDTH-1:0] out131,
  output [WIDTH-1:0] out132,
  output [WIDTH-1:0] out133,
  output [WIDTH-1:0] out134,
  output [WIDTH-1:0] out135,
  output [WIDTH-1:0] out136,
  output [WIDTH-1:0] out137,
  output [WIDTH-1:0] out138,
  output [WIDTH-1:0] out139,
  output [WIDTH-1:0] out140,
  output [WIDTH-1:0] out141,
  output [WIDTH-1:0] out142,
  output [WIDTH-1:0] out143,
  output [WIDTH-1:0] out144,
  output [WIDTH-1:0] out145,
  output [WIDTH-1:0] out146,
  output [WIDTH-1:0] out147,
  output [WIDTH-1:0] out148,
  output [WIDTH-1:0] out149,
  output [WIDTH-1:0] out150,
  output [WIDTH-1:0] out151,
  output [WIDTH-1:0] out152,
  output [WIDTH-1:0] out153,
  output [WIDTH-1:0] out154,
  output [WIDTH-1:0] out155,
  output [WIDTH-1:0] out156,
  output [WIDTH-1:0] out157,
  output [WIDTH-1:0] out158,
  output [WIDTH-1:0] out159,
  output [WIDTH-1:0] out160,
  output [WIDTH-1:0] out161,
  output [WIDTH-1:0] out162,
  output [WIDTH-1:0] out163,
  output [WIDTH-1:0] out164,
  output [WIDTH-1:0] out165,
  output [WIDTH-1:0] out166,
  output [WIDTH-1:0] out167,
  output [WIDTH-1:0] out168,
  output [WIDTH-1:0] out169,
  output [WIDTH-1:0] out170,
  output [WIDTH-1:0] out171,
  output [WIDTH-1:0] out172,
  output [WIDTH-1:0] out173,
  output [WIDTH-1:0] out174,
  output [WIDTH-1:0] out175,
  output [WIDTH-1:0] out176,
  output [WIDTH-1:0] out177,
  output [WIDTH-1:0] out178,
  output [WIDTH-1:0] out179,
  output [WIDTH-1:0] out180,
  output [WIDTH-1:0] out181,
  output [WIDTH-1:0] out182,
  output [WIDTH-1:0] out183,
  output [WIDTH-1:0] out184,
  output [WIDTH-1:0] out185,
  output [WIDTH-1:0] out186,
  output [WIDTH-1:0] out187,
  output [WIDTH-1:0] out188,
  output [WIDTH-1:0] out189,
  output [WIDTH-1:0] out190,
  output [WIDTH-1:0] out191,
  output [WIDTH-1:0] out192,
  output [WIDTH-1:0] out193,
  output [WIDTH-1:0] out194,
  output [WIDTH-1:0] out195,
  output [WIDTH-1:0] out196,
  output [WIDTH-1:0] out197,
  output [WIDTH-1:0] out198,
  output [WIDTH-1:0] out199,
  output [WIDTH-1:0] out200,
  output [WIDTH-1:0] out201,
  output [WIDTH-1:0] out202,
  output [WIDTH-1:0] out203,
  output [WIDTH-1:0] out204,
  output [WIDTH-1:0] out205,
  output [WIDTH-1:0] out206,
  output [WIDTH-1:0] out207,
  output [WIDTH-1:0] out208,
  output [WIDTH-1:0] out209,
  output [WIDTH-1:0] out210,
  output [WIDTH-1:0] out211,
  output [WIDTH-1:0] out212,
  output [WIDTH-1:0] out213,
  output [WIDTH-1:0] out214,
  output [WIDTH-1:0] out215,
  output [WIDTH-1:0] out216,
  output [WIDTH-1:0] out217,
  output [WIDTH-1:0] out218,
  output [WIDTH-1:0] out219,
  output [WIDTH-1:0] out220,
  output [WIDTH-1:0] out221,
  output [WIDTH-1:0] out222,
  output [WIDTH-1:0] out223,
  output [WIDTH-1:0] out224,
  output [WIDTH-1:0] out225,
  output [WIDTH-1:0] out226,
  output [WIDTH-1:0] out227,
  output [WIDTH-1:0] out228,
  output [WIDTH-1:0] out229,
  output [WIDTH-1:0] out230,
  output [WIDTH-1:0] out231,
  output [WIDTH-1:0] out232,
  output [WIDTH-1:0] out233,
  output [WIDTH-1:0] out234,
  output [WIDTH-1:0] out235,
  output [WIDTH-1:0] out236,
  output [WIDTH-1:0] out237,
  output [WIDTH-1:0] out238,
  output [WIDTH-1:0] out239,
  output [WIDTH-1:0] out240,
  output [WIDTH-1:0] out241,
  output [WIDTH-1:0] out242,
  output [WIDTH-1:0] out243,
  output [WIDTH-1:0] out244,
  output [WIDTH-1:0] out245,
  output [WIDTH-1:0] out246,
  output [WIDTH-1:0] out247,
  output [WIDTH-1:0] out248,
  output [WIDTH-1:0] out249,
  output [WIDTH-1:0] out250,
  output [WIDTH-1:0] out251,
  output [WIDTH-1:0] out252,
  output [WIDTH-1:0] out253,
  output [WIDTH-1:0] out254,
  output [WIDTH-1:0] out255
);

  wire [2304-1:0] conf_out;
  wire [WIDTH-1:0] in_reg_wire_0 [0:256-1];
  wire [WIDTH-1:0] in_reg_wire_1 [0:256-1];
  wire [WIDTH-1:0] in_reg_wire_2 [0:256-1];
  wire [WIDTH-1:0] in_reg_wire_3 [0:256-1];
  wire [WIDTH-1:0] in_reg_wire_4 [0:256-1];
  wire [WIDTH-1:0] in_reg_wire_5 [0:256-1];
  wire [64-1:0] net_conf_bus [0:96-1];

  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg0
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus_in),
    .out(net_conf_bus[0])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(1),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_0
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[0]),
    .swicth_conf_out(conf_out[23:0])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg1
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[0]),
    .out(net_conf_bus[1])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(2),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_1
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[1]),
    .swicth_conf_out(conf_out[47:24])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg2
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[1]),
    .out(net_conf_bus[2])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(3),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_2
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[2]),
    .swicth_conf_out(conf_out[71:48])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg3
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[2]),
    .out(net_conf_bus[3])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(4),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_3
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[3]),
    .swicth_conf_out(conf_out[95:72])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg4
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[3]),
    .out(net_conf_bus[4])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(5),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_4
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[4]),
    .swicth_conf_out(conf_out[119:96])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg5
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[4]),
    .out(net_conf_bus[5])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(6),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_5
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[5]),
    .swicth_conf_out(conf_out[143:120])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg6
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[5]),
    .out(net_conf_bus[6])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(7),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_6
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[6]),
    .swicth_conf_out(conf_out[167:144])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg7
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[6]),
    .out(net_conf_bus[7])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(8),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_7
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[7]),
    .swicth_conf_out(conf_out[191:168])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg8
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[7]),
    .out(net_conf_bus[8])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(9),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_8
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[8]),
    .swicth_conf_out(conf_out[215:192])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg9
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[8]),
    .out(net_conf_bus[9])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(10),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_9
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[9]),
    .swicth_conf_out(conf_out[239:216])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg10
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[9]),
    .out(net_conf_bus[10])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(11),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_10
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[10]),
    .swicth_conf_out(conf_out[263:240])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg11
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[10]),
    .out(net_conf_bus[11])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(12),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_11
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[11]),
    .swicth_conf_out(conf_out[287:264])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg12
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[11]),
    .out(net_conf_bus[12])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(13),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_12
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[12]),
    .swicth_conf_out(conf_out[311:288])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg13
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[12]),
    .out(net_conf_bus[13])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(14),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_13
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[13]),
    .swicth_conf_out(conf_out[335:312])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg14
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[13]),
    .out(net_conf_bus[14])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(15),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_14
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[14]),
    .swicth_conf_out(conf_out[359:336])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg15
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[14]),
    .out(net_conf_bus[15])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(16),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_15
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[15]),
    .swicth_conf_out(conf_out[383:360])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg16
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[15]),
    .out(net_conf_bus[16])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(17),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_16
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[16]),
    .swicth_conf_out(conf_out[407:384])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg17
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[16]),
    .out(net_conf_bus[17])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(18),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_17
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[17]),
    .swicth_conf_out(conf_out[431:408])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg18
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[17]),
    .out(net_conf_bus[18])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(19),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_18
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[18]),
    .swicth_conf_out(conf_out[455:432])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg19
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[18]),
    .out(net_conf_bus[19])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(20),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_19
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[19]),
    .swicth_conf_out(conf_out[479:456])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg20
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[19]),
    .out(net_conf_bus[20])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(21),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_20
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[20]),
    .swicth_conf_out(conf_out[503:480])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg21
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[20]),
    .out(net_conf_bus[21])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(22),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_21
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[21]),
    .swicth_conf_out(conf_out[527:504])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg22
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[21]),
    .out(net_conf_bus[22])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(23),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_22
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[22]),
    .swicth_conf_out(conf_out[551:528])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg23
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[22]),
    .out(net_conf_bus[23])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(24),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_23
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[23]),
    .swicth_conf_out(conf_out[575:552])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg24
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[23]),
    .out(net_conf_bus[24])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(25),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_24
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[24]),
    .swicth_conf_out(conf_out[599:576])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg25
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[24]),
    .out(net_conf_bus[25])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(26),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_25
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[25]),
    .swicth_conf_out(conf_out[623:600])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg26
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[25]),
    .out(net_conf_bus[26])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(27),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_26
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[26]),
    .swicth_conf_out(conf_out[647:624])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg27
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[26]),
    .out(net_conf_bus[27])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(28),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_27
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[27]),
    .swicth_conf_out(conf_out[671:648])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg28
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[27]),
    .out(net_conf_bus[28])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(29),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_28
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[28]),
    .swicth_conf_out(conf_out[695:672])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg29
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[28]),
    .out(net_conf_bus[29])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(30),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_29
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[29]),
    .swicth_conf_out(conf_out[719:696])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg30
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[29]),
    .out(net_conf_bus[30])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(31),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_30
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[30]),
    .swicth_conf_out(conf_out[743:720])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg31
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[30]),
    .out(net_conf_bus[31])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(32),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_31
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[31]),
    .swicth_conf_out(conf_out[767:744])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg32
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[31]),
    .out(net_conf_bus[32])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(33),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_32
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[32]),
    .swicth_conf_out(conf_out[791:768])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg33
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[32]),
    .out(net_conf_bus[33])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(34),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_33
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[33]),
    .swicth_conf_out(conf_out[815:792])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg34
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[33]),
    .out(net_conf_bus[34])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(35),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_34
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[34]),
    .swicth_conf_out(conf_out[839:816])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg35
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[34]),
    .out(net_conf_bus[35])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(36),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_35
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[35]),
    .swicth_conf_out(conf_out[863:840])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg36
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[35]),
    .out(net_conf_bus[36])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(37),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_36
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[36]),
    .swicth_conf_out(conf_out[887:864])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg37
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[36]),
    .out(net_conf_bus[37])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(38),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_37
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[37]),
    .swicth_conf_out(conf_out[911:888])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg38
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[37]),
    .out(net_conf_bus[38])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(39),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_38
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[38]),
    .swicth_conf_out(conf_out[935:912])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg39
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[38]),
    .out(net_conf_bus[39])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(40),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_39
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[39]),
    .swicth_conf_out(conf_out[959:936])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg40
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[39]),
    .out(net_conf_bus[40])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(41),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_40
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[40]),
    .swicth_conf_out(conf_out[983:960])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg41
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[40]),
    .out(net_conf_bus[41])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(42),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_41
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[41]),
    .swicth_conf_out(conf_out[1007:984])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg42
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[41]),
    .out(net_conf_bus[42])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(43),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_42
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[42]),
    .swicth_conf_out(conf_out[1031:1008])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg43
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[42]),
    .out(net_conf_bus[43])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(44),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_43
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[43]),
    .swicth_conf_out(conf_out[1055:1032])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg44
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[43]),
    .out(net_conf_bus[44])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(45),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_44
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[44]),
    .swicth_conf_out(conf_out[1079:1056])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg45
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[44]),
    .out(net_conf_bus[45])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(46),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_45
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[45]),
    .swicth_conf_out(conf_out[1103:1080])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg46
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[45]),
    .out(net_conf_bus[46])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(47),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_46
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[46]),
    .swicth_conf_out(conf_out[1127:1104])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg47
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[46]),
    .out(net_conf_bus[47])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(48),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_47
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[47]),
    .swicth_conf_out(conf_out[1151:1128])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg48
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[47]),
    .out(net_conf_bus[48])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(49),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_48
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[48]),
    .swicth_conf_out(conf_out[1175:1152])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg49
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[48]),
    .out(net_conf_bus[49])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(50),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_49
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[49]),
    .swicth_conf_out(conf_out[1199:1176])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg50
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[49]),
    .out(net_conf_bus[50])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(51),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_50
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[50]),
    .swicth_conf_out(conf_out[1223:1200])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg51
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[50]),
    .out(net_conf_bus[51])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(52),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_51
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[51]),
    .swicth_conf_out(conf_out[1247:1224])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg52
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[51]),
    .out(net_conf_bus[52])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(53),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_52
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[52]),
    .swicth_conf_out(conf_out[1271:1248])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg53
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[52]),
    .out(net_conf_bus[53])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(54),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_53
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[53]),
    .swicth_conf_out(conf_out[1295:1272])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg54
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[53]),
    .out(net_conf_bus[54])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(55),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_54
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[54]),
    .swicth_conf_out(conf_out[1319:1296])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg55
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[54]),
    .out(net_conf_bus[55])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(56),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_55
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[55]),
    .swicth_conf_out(conf_out[1343:1320])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg56
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[55]),
    .out(net_conf_bus[56])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(57),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_56
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[56]),
    .swicth_conf_out(conf_out[1367:1344])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg57
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[56]),
    .out(net_conf_bus[57])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(58),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_57
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[57]),
    .swicth_conf_out(conf_out[1391:1368])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg58
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[57]),
    .out(net_conf_bus[58])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(59),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_58
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[58]),
    .swicth_conf_out(conf_out[1415:1392])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg59
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[58]),
    .out(net_conf_bus[59])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(60),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_59
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[59]),
    .swicth_conf_out(conf_out[1439:1416])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg60
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[59]),
    .out(net_conf_bus[60])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(61),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_60
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[60]),
    .swicth_conf_out(conf_out[1463:1440])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg61
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[60]),
    .out(net_conf_bus[61])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(62),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_61
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[61]),
    .swicth_conf_out(conf_out[1487:1464])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg62
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[61]),
    .out(net_conf_bus[62])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(63),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_62
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[62]),
    .swicth_conf_out(conf_out[1511:1488])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg63
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[62]),
    .out(net_conf_bus[63])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(64),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_63
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[63]),
    .swicth_conf_out(conf_out[1535:1512])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg64
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[63]),
    .out(net_conf_bus[64])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(65),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_64
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[64]),
    .swicth_conf_out(conf_out[1559:1536])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg65
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[64]),
    .out(net_conf_bus[65])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(66),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_65
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[65]),
    .swicth_conf_out(conf_out[1583:1560])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg66
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[65]),
    .out(net_conf_bus[66])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(67),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_66
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[66]),
    .swicth_conf_out(conf_out[1607:1584])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg67
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[66]),
    .out(net_conf_bus[67])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(68),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_67
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[67]),
    .swicth_conf_out(conf_out[1631:1608])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg68
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[67]),
    .out(net_conf_bus[68])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(69),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_68
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[68]),
    .swicth_conf_out(conf_out[1655:1632])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg69
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[68]),
    .out(net_conf_bus[69])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(70),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_69
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[69]),
    .swicth_conf_out(conf_out[1679:1656])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg70
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[69]),
    .out(net_conf_bus[70])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(71),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_70
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[70]),
    .swicth_conf_out(conf_out[1703:1680])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg71
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[70]),
    .out(net_conf_bus[71])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(72),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_71
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[71]),
    .swicth_conf_out(conf_out[1727:1704])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg72
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[71]),
    .out(net_conf_bus[72])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(73),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_72
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[72]),
    .swicth_conf_out(conf_out[1751:1728])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg73
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[72]),
    .out(net_conf_bus[73])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(74),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_73
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[73]),
    .swicth_conf_out(conf_out[1775:1752])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg74
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[73]),
    .out(net_conf_bus[74])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(75),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_74
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[74]),
    .swicth_conf_out(conf_out[1799:1776])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg75
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[74]),
    .out(net_conf_bus[75])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(76),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_75
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[75]),
    .swicth_conf_out(conf_out[1823:1800])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg76
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[75]),
    .out(net_conf_bus[76])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(77),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_76
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[76]),
    .swicth_conf_out(conf_out[1847:1824])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg77
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[76]),
    .out(net_conf_bus[77])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(78),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_77
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[77]),
    .swicth_conf_out(conf_out[1871:1848])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg78
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[77]),
    .out(net_conf_bus[78])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(79),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_78
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[78]),
    .swicth_conf_out(conf_out[1895:1872])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg79
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[78]),
    .out(net_conf_bus[79])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(80),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_79
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[79]),
    .swicth_conf_out(conf_out[1919:1896])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg80
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[79]),
    .out(net_conf_bus[80])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(81),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_80
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[80]),
    .swicth_conf_out(conf_out[1943:1920])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg81
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[80]),
    .out(net_conf_bus[81])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(82),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_81
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[81]),
    .swicth_conf_out(conf_out[1967:1944])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg82
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[81]),
    .out(net_conf_bus[82])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(83),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_82
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[82]),
    .swicth_conf_out(conf_out[1991:1968])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg83
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[82]),
    .out(net_conf_bus[83])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(84),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_83
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[83]),
    .swicth_conf_out(conf_out[2015:1992])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg84
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[83]),
    .out(net_conf_bus[84])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(85),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_84
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[84]),
    .swicth_conf_out(conf_out[2039:2016])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg85
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[84]),
    .out(net_conf_bus[85])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(86),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_85
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[85]),
    .swicth_conf_out(conf_out[2063:2040])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg86
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[85]),
    .out(net_conf_bus[86])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(87),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_86
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[86]),
    .swicth_conf_out(conf_out[2087:2064])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg87
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[86]),
    .out(net_conf_bus[87])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(88),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_87
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[87]),
    .swicth_conf_out(conf_out[2111:2088])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg88
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[87]),
    .out(net_conf_bus[88])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(89),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_88
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[88]),
    .swicth_conf_out(conf_out[2135:2112])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg89
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[88]),
    .out(net_conf_bus[89])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(90),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_89
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[89]),
    .swicth_conf_out(conf_out[2159:2136])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg90
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[89]),
    .out(net_conf_bus[90])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(91),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_90
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[90]),
    .swicth_conf_out(conf_out[2183:2160])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg91
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[90]),
    .out(net_conf_bus[91])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(92),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_91
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[91]),
    .swicth_conf_out(conf_out[2207:2184])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg92
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[91]),
    .out(net_conf_bus[92])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(93),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_92
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[92]),
    .swicth_conf_out(conf_out[2231:2208])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg93
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[92]),
    .out(net_conf_bus[93])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(94),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_93
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[93]),
    .swicth_conf_out(conf_out[2255:2232])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg94
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[93]),
    .out(net_conf_bus[94])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(95),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_94
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[94]),
    .swicth_conf_out(conf_out[2279:2256])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg95
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[94]),
    .out(net_conf_bus[95])
  );


  swicth_conf_control_24_1
  #(
    .SWICTH_NUMBER(96),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_95
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[95]),
    .swicth_conf_out(conf_out[2303:2280])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_0
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in0),
    .out(in_reg_wire_0[0])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_1
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in1),
    .out(in_reg_wire_0[1])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_2
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in2),
    .out(in_reg_wire_0[2])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_3
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in3),
    .out(in_reg_wire_0[3])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_4
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in4),
    .out(in_reg_wire_0[4])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_5
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in5),
    .out(in_reg_wire_0[5])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_6
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in6),
    .out(in_reg_wire_0[6])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_7
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in7),
    .out(in_reg_wire_0[7])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_8
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in8),
    .out(in_reg_wire_0[8])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_9
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in9),
    .out(in_reg_wire_0[9])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_10
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in10),
    .out(in_reg_wire_0[10])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_11
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in11),
    .out(in_reg_wire_0[11])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_12
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in12),
    .out(in_reg_wire_0[12])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_13
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in13),
    .out(in_reg_wire_0[13])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_14
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in14),
    .out(in_reg_wire_0[14])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_15
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in15),
    .out(in_reg_wire_0[15])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_16
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in16),
    .out(in_reg_wire_0[16])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_17
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in17),
    .out(in_reg_wire_0[17])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_18
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in18),
    .out(in_reg_wire_0[18])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_19
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in19),
    .out(in_reg_wire_0[19])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_20
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in20),
    .out(in_reg_wire_0[20])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_21
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in21),
    .out(in_reg_wire_0[21])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_22
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in22),
    .out(in_reg_wire_0[22])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_23
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in23),
    .out(in_reg_wire_0[23])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_24
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in24),
    .out(in_reg_wire_0[24])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_25
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in25),
    .out(in_reg_wire_0[25])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_26
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in26),
    .out(in_reg_wire_0[26])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_27
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in27),
    .out(in_reg_wire_0[27])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_28
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in28),
    .out(in_reg_wire_0[28])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_29
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in29),
    .out(in_reg_wire_0[29])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_30
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in30),
    .out(in_reg_wire_0[30])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_31
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in31),
    .out(in_reg_wire_0[31])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_32
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in32),
    .out(in_reg_wire_0[32])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_33
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in33),
    .out(in_reg_wire_0[33])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_34
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in34),
    .out(in_reg_wire_0[34])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_35
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in35),
    .out(in_reg_wire_0[35])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_36
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in36),
    .out(in_reg_wire_0[36])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_37
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in37),
    .out(in_reg_wire_0[37])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_38
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in38),
    .out(in_reg_wire_0[38])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_39
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in39),
    .out(in_reg_wire_0[39])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_40
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in40),
    .out(in_reg_wire_0[40])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_41
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in41),
    .out(in_reg_wire_0[41])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_42
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in42),
    .out(in_reg_wire_0[42])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_43
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in43),
    .out(in_reg_wire_0[43])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_44
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in44),
    .out(in_reg_wire_0[44])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_45
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in45),
    .out(in_reg_wire_0[45])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_46
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in46),
    .out(in_reg_wire_0[46])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_47
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in47),
    .out(in_reg_wire_0[47])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_48
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in48),
    .out(in_reg_wire_0[48])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_49
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in49),
    .out(in_reg_wire_0[49])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_50
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in50),
    .out(in_reg_wire_0[50])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_51
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in51),
    .out(in_reg_wire_0[51])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_52
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in52),
    .out(in_reg_wire_0[52])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_53
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in53),
    .out(in_reg_wire_0[53])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_54
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in54),
    .out(in_reg_wire_0[54])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_55
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in55),
    .out(in_reg_wire_0[55])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_56
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in56),
    .out(in_reg_wire_0[56])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_57
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in57),
    .out(in_reg_wire_0[57])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_58
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in58),
    .out(in_reg_wire_0[58])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_59
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in59),
    .out(in_reg_wire_0[59])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_60
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in60),
    .out(in_reg_wire_0[60])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_61
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in61),
    .out(in_reg_wire_0[61])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_62
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in62),
    .out(in_reg_wire_0[62])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_63
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in63),
    .out(in_reg_wire_0[63])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_64
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in64),
    .out(in_reg_wire_0[64])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_65
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in65),
    .out(in_reg_wire_0[65])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_66
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in66),
    .out(in_reg_wire_0[66])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_67
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in67),
    .out(in_reg_wire_0[67])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_68
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in68),
    .out(in_reg_wire_0[68])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_69
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in69),
    .out(in_reg_wire_0[69])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_70
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in70),
    .out(in_reg_wire_0[70])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_71
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in71),
    .out(in_reg_wire_0[71])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_72
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in72),
    .out(in_reg_wire_0[72])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_73
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in73),
    .out(in_reg_wire_0[73])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_74
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in74),
    .out(in_reg_wire_0[74])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_75
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in75),
    .out(in_reg_wire_0[75])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_76
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in76),
    .out(in_reg_wire_0[76])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_77
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in77),
    .out(in_reg_wire_0[77])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_78
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in78),
    .out(in_reg_wire_0[78])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_79
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in79),
    .out(in_reg_wire_0[79])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_80
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in80),
    .out(in_reg_wire_0[80])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_81
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in81),
    .out(in_reg_wire_0[81])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_82
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in82),
    .out(in_reg_wire_0[82])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_83
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in83),
    .out(in_reg_wire_0[83])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_84
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in84),
    .out(in_reg_wire_0[84])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_85
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in85),
    .out(in_reg_wire_0[85])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_86
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in86),
    .out(in_reg_wire_0[86])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_87
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in87),
    .out(in_reg_wire_0[87])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_88
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in88),
    .out(in_reg_wire_0[88])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_89
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in89),
    .out(in_reg_wire_0[89])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_90
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in90),
    .out(in_reg_wire_0[90])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_91
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in91),
    .out(in_reg_wire_0[91])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_92
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in92),
    .out(in_reg_wire_0[92])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_93
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in93),
    .out(in_reg_wire_0[93])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_94
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in94),
    .out(in_reg_wire_0[94])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_95
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in95),
    .out(in_reg_wire_0[95])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_96
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in96),
    .out(in_reg_wire_0[96])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_97
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in97),
    .out(in_reg_wire_0[97])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_98
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in98),
    .out(in_reg_wire_0[98])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_99
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in99),
    .out(in_reg_wire_0[99])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_100
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in100),
    .out(in_reg_wire_0[100])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_101
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in101),
    .out(in_reg_wire_0[101])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_102
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in102),
    .out(in_reg_wire_0[102])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_103
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in103),
    .out(in_reg_wire_0[103])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_104
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in104),
    .out(in_reg_wire_0[104])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_105
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in105),
    .out(in_reg_wire_0[105])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_106
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in106),
    .out(in_reg_wire_0[106])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_107
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in107),
    .out(in_reg_wire_0[107])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_108
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in108),
    .out(in_reg_wire_0[108])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_109
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in109),
    .out(in_reg_wire_0[109])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_110
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in110),
    .out(in_reg_wire_0[110])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_111
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in111),
    .out(in_reg_wire_0[111])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_112
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in112),
    .out(in_reg_wire_0[112])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_113
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in113),
    .out(in_reg_wire_0[113])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_114
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in114),
    .out(in_reg_wire_0[114])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_115
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in115),
    .out(in_reg_wire_0[115])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_116
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in116),
    .out(in_reg_wire_0[116])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_117
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in117),
    .out(in_reg_wire_0[117])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_118
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in118),
    .out(in_reg_wire_0[118])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_119
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in119),
    .out(in_reg_wire_0[119])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_120
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in120),
    .out(in_reg_wire_0[120])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_121
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in121),
    .out(in_reg_wire_0[121])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_122
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in122),
    .out(in_reg_wire_0[122])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_123
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in123),
    .out(in_reg_wire_0[123])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_124
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in124),
    .out(in_reg_wire_0[124])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_125
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in125),
    .out(in_reg_wire_0[125])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_126
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in126),
    .out(in_reg_wire_0[126])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_127
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in127),
    .out(in_reg_wire_0[127])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_128
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in128),
    .out(in_reg_wire_0[128])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_129
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in129),
    .out(in_reg_wire_0[129])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_130
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in130),
    .out(in_reg_wire_0[130])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_131
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in131),
    .out(in_reg_wire_0[131])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_132
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in132),
    .out(in_reg_wire_0[132])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_133
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in133),
    .out(in_reg_wire_0[133])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_134
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in134),
    .out(in_reg_wire_0[134])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_135
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in135),
    .out(in_reg_wire_0[135])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_136
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in136),
    .out(in_reg_wire_0[136])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_137
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in137),
    .out(in_reg_wire_0[137])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_138
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in138),
    .out(in_reg_wire_0[138])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_139
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in139),
    .out(in_reg_wire_0[139])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_140
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in140),
    .out(in_reg_wire_0[140])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_141
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in141),
    .out(in_reg_wire_0[141])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_142
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in142),
    .out(in_reg_wire_0[142])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_143
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in143),
    .out(in_reg_wire_0[143])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_144
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in144),
    .out(in_reg_wire_0[144])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_145
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in145),
    .out(in_reg_wire_0[145])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_146
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in146),
    .out(in_reg_wire_0[146])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_147
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in147),
    .out(in_reg_wire_0[147])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_148
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in148),
    .out(in_reg_wire_0[148])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_149
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in149),
    .out(in_reg_wire_0[149])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_150
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in150),
    .out(in_reg_wire_0[150])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_151
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in151),
    .out(in_reg_wire_0[151])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_152
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in152),
    .out(in_reg_wire_0[152])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_153
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in153),
    .out(in_reg_wire_0[153])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_154
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in154),
    .out(in_reg_wire_0[154])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_155
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in155),
    .out(in_reg_wire_0[155])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_156
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in156),
    .out(in_reg_wire_0[156])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_157
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in157),
    .out(in_reg_wire_0[157])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_158
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in158),
    .out(in_reg_wire_0[158])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_159
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in159),
    .out(in_reg_wire_0[159])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_160
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in160),
    .out(in_reg_wire_0[160])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_161
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in161),
    .out(in_reg_wire_0[161])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_162
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in162),
    .out(in_reg_wire_0[162])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_163
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in163),
    .out(in_reg_wire_0[163])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_164
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in164),
    .out(in_reg_wire_0[164])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_165
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in165),
    .out(in_reg_wire_0[165])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_166
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in166),
    .out(in_reg_wire_0[166])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_167
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in167),
    .out(in_reg_wire_0[167])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_168
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in168),
    .out(in_reg_wire_0[168])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_169
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in169),
    .out(in_reg_wire_0[169])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_170
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in170),
    .out(in_reg_wire_0[170])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_171
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in171),
    .out(in_reg_wire_0[171])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_172
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in172),
    .out(in_reg_wire_0[172])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_173
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in173),
    .out(in_reg_wire_0[173])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_174
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in174),
    .out(in_reg_wire_0[174])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_175
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in175),
    .out(in_reg_wire_0[175])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_176
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in176),
    .out(in_reg_wire_0[176])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_177
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in177),
    .out(in_reg_wire_0[177])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_178
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in178),
    .out(in_reg_wire_0[178])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_179
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in179),
    .out(in_reg_wire_0[179])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_180
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in180),
    .out(in_reg_wire_0[180])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_181
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in181),
    .out(in_reg_wire_0[181])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_182
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in182),
    .out(in_reg_wire_0[182])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_183
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in183),
    .out(in_reg_wire_0[183])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_184
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in184),
    .out(in_reg_wire_0[184])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_185
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in185),
    .out(in_reg_wire_0[185])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_186
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in186),
    .out(in_reg_wire_0[186])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_187
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in187),
    .out(in_reg_wire_0[187])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_188
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in188),
    .out(in_reg_wire_0[188])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_189
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in189),
    .out(in_reg_wire_0[189])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_190
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in190),
    .out(in_reg_wire_0[190])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_191
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in191),
    .out(in_reg_wire_0[191])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_192
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in192),
    .out(in_reg_wire_0[192])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_193
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in193),
    .out(in_reg_wire_0[193])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_194
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in194),
    .out(in_reg_wire_0[194])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_195
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in195),
    .out(in_reg_wire_0[195])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_196
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in196),
    .out(in_reg_wire_0[196])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_197
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in197),
    .out(in_reg_wire_0[197])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_198
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in198),
    .out(in_reg_wire_0[198])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_199
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in199),
    .out(in_reg_wire_0[199])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_200
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in200),
    .out(in_reg_wire_0[200])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_201
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in201),
    .out(in_reg_wire_0[201])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_202
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in202),
    .out(in_reg_wire_0[202])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_203
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in203),
    .out(in_reg_wire_0[203])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_204
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in204),
    .out(in_reg_wire_0[204])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_205
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in205),
    .out(in_reg_wire_0[205])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_206
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in206),
    .out(in_reg_wire_0[206])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_207
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in207),
    .out(in_reg_wire_0[207])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_208
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in208),
    .out(in_reg_wire_0[208])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_209
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in209),
    .out(in_reg_wire_0[209])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_210
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in210),
    .out(in_reg_wire_0[210])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_211
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in211),
    .out(in_reg_wire_0[211])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_212
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in212),
    .out(in_reg_wire_0[212])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_213
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in213),
    .out(in_reg_wire_0[213])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_214
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in214),
    .out(in_reg_wire_0[214])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_215
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in215),
    .out(in_reg_wire_0[215])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_216
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in216),
    .out(in_reg_wire_0[216])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_217
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in217),
    .out(in_reg_wire_0[217])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_218
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in218),
    .out(in_reg_wire_0[218])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_219
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in219),
    .out(in_reg_wire_0[219])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_220
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in220),
    .out(in_reg_wire_0[220])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_221
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in221),
    .out(in_reg_wire_0[221])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_222
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in222),
    .out(in_reg_wire_0[222])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_223
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in223),
    .out(in_reg_wire_0[223])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_224
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in224),
    .out(in_reg_wire_0[224])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_225
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in225),
    .out(in_reg_wire_0[225])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_226
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in226),
    .out(in_reg_wire_0[226])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_227
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in227),
    .out(in_reg_wire_0[227])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_228
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in228),
    .out(in_reg_wire_0[228])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_229
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in229),
    .out(in_reg_wire_0[229])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_230
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in230),
    .out(in_reg_wire_0[230])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_231
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in231),
    .out(in_reg_wire_0[231])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_232
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in232),
    .out(in_reg_wire_0[232])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_233
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in233),
    .out(in_reg_wire_0[233])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_234
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in234),
    .out(in_reg_wire_0[234])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_235
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in235),
    .out(in_reg_wire_0[235])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_236
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in236),
    .out(in_reg_wire_0[236])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_237
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in237),
    .out(in_reg_wire_0[237])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_238
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in238),
    .out(in_reg_wire_0[238])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_239
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in239),
    .out(in_reg_wire_0[239])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_240
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in240),
    .out(in_reg_wire_0[240])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_241
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in241),
    .out(in_reg_wire_0[241])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_242
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in242),
    .out(in_reg_wire_0[242])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_243
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in243),
    .out(in_reg_wire_0[243])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_244
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in244),
    .out(in_reg_wire_0[244])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_245
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in245),
    .out(in_reg_wire_0[245])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_246
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in246),
    .out(in_reg_wire_0[246])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_247
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in247),
    .out(in_reg_wire_0[247])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_248
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in248),
    .out(in_reg_wire_0[248])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_249
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in249),
    .out(in_reg_wire_0[249])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_250
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in250),
    .out(in_reg_wire_0[250])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_251
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in251),
    .out(in_reg_wire_0[251])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_252
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in252),
    .out(in_reg_wire_0[252])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_253
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in253),
    .out(in_reg_wire_0[253])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_254
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in254),
    .out(in_reg_wire_0[254])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_255
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in255),
    .out(in_reg_wire_0[255])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_0
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[0]),
    .out(in_reg_wire_2[0])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_1
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[1]),
    .out(in_reg_wire_2[1])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_2
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[2]),
    .out(in_reg_wire_2[2])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_3
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[3]),
    .out(in_reg_wire_2[3])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_4
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[4]),
    .out(in_reg_wire_2[4])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_5
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[5]),
    .out(in_reg_wire_2[5])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_6
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[6]),
    .out(in_reg_wire_2[6])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_7
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[7]),
    .out(in_reg_wire_2[7])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_8
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[8]),
    .out(in_reg_wire_2[8])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_9
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[9]),
    .out(in_reg_wire_2[9])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_10
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[10]),
    .out(in_reg_wire_2[10])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_11
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[11]),
    .out(in_reg_wire_2[11])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_12
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[12]),
    .out(in_reg_wire_2[12])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_13
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[13]),
    .out(in_reg_wire_2[13])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_14
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[14]),
    .out(in_reg_wire_2[14])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_15
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[15]),
    .out(in_reg_wire_2[15])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_16
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[16]),
    .out(in_reg_wire_2[16])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_17
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[17]),
    .out(in_reg_wire_2[17])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_18
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[18]),
    .out(in_reg_wire_2[18])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_19
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[19]),
    .out(in_reg_wire_2[19])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_20
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[20]),
    .out(in_reg_wire_2[20])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_21
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[21]),
    .out(in_reg_wire_2[21])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_22
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[22]),
    .out(in_reg_wire_2[22])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_23
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[23]),
    .out(in_reg_wire_2[23])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_24
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[24]),
    .out(in_reg_wire_2[24])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_25
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[25]),
    .out(in_reg_wire_2[25])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_26
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[26]),
    .out(in_reg_wire_2[26])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_27
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[27]),
    .out(in_reg_wire_2[27])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_28
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[28]),
    .out(in_reg_wire_2[28])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_29
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[29]),
    .out(in_reg_wire_2[29])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_30
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[30]),
    .out(in_reg_wire_2[30])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_31
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[31]),
    .out(in_reg_wire_2[31])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_32
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[32]),
    .out(in_reg_wire_2[32])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_33
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[33]),
    .out(in_reg_wire_2[33])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_34
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[34]),
    .out(in_reg_wire_2[34])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_35
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[35]),
    .out(in_reg_wire_2[35])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_36
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[36]),
    .out(in_reg_wire_2[36])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_37
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[37]),
    .out(in_reg_wire_2[37])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_38
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[38]),
    .out(in_reg_wire_2[38])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_39
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[39]),
    .out(in_reg_wire_2[39])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_40
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[40]),
    .out(in_reg_wire_2[40])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_41
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[41]),
    .out(in_reg_wire_2[41])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_42
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[42]),
    .out(in_reg_wire_2[42])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_43
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[43]),
    .out(in_reg_wire_2[43])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_44
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[44]),
    .out(in_reg_wire_2[44])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_45
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[45]),
    .out(in_reg_wire_2[45])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_46
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[46]),
    .out(in_reg_wire_2[46])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_47
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[47]),
    .out(in_reg_wire_2[47])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_48
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[48]),
    .out(in_reg_wire_2[48])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_49
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[49]),
    .out(in_reg_wire_2[49])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_50
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[50]),
    .out(in_reg_wire_2[50])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_51
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[51]),
    .out(in_reg_wire_2[51])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_52
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[52]),
    .out(in_reg_wire_2[52])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_53
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[53]),
    .out(in_reg_wire_2[53])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_54
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[54]),
    .out(in_reg_wire_2[54])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_55
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[55]),
    .out(in_reg_wire_2[55])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_56
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[56]),
    .out(in_reg_wire_2[56])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_57
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[57]),
    .out(in_reg_wire_2[57])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_58
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[58]),
    .out(in_reg_wire_2[58])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_59
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[59]),
    .out(in_reg_wire_2[59])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_60
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[60]),
    .out(in_reg_wire_2[60])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_61
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[61]),
    .out(in_reg_wire_2[61])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_62
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[62]),
    .out(in_reg_wire_2[62])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_63
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[63]),
    .out(in_reg_wire_2[63])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_64
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[64]),
    .out(in_reg_wire_2[64])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_65
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[65]),
    .out(in_reg_wire_2[65])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_66
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[66]),
    .out(in_reg_wire_2[66])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_67
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[67]),
    .out(in_reg_wire_2[67])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_68
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[68]),
    .out(in_reg_wire_2[68])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_69
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[69]),
    .out(in_reg_wire_2[69])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_70
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[70]),
    .out(in_reg_wire_2[70])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_71
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[71]),
    .out(in_reg_wire_2[71])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_72
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[72]),
    .out(in_reg_wire_2[72])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_73
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[73]),
    .out(in_reg_wire_2[73])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_74
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[74]),
    .out(in_reg_wire_2[74])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_75
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[75]),
    .out(in_reg_wire_2[75])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_76
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[76]),
    .out(in_reg_wire_2[76])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_77
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[77]),
    .out(in_reg_wire_2[77])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_78
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[78]),
    .out(in_reg_wire_2[78])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_79
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[79]),
    .out(in_reg_wire_2[79])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_80
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[80]),
    .out(in_reg_wire_2[80])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_81
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[81]),
    .out(in_reg_wire_2[81])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_82
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[82]),
    .out(in_reg_wire_2[82])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_83
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[83]),
    .out(in_reg_wire_2[83])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_84
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[84]),
    .out(in_reg_wire_2[84])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_85
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[85]),
    .out(in_reg_wire_2[85])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_86
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[86]),
    .out(in_reg_wire_2[86])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_87
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[87]),
    .out(in_reg_wire_2[87])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_88
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[88]),
    .out(in_reg_wire_2[88])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_89
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[89]),
    .out(in_reg_wire_2[89])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_90
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[90]),
    .out(in_reg_wire_2[90])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_91
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[91]),
    .out(in_reg_wire_2[91])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_92
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[92]),
    .out(in_reg_wire_2[92])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_93
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[93]),
    .out(in_reg_wire_2[93])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_94
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[94]),
    .out(in_reg_wire_2[94])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_95
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[95]),
    .out(in_reg_wire_2[95])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_96
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[96]),
    .out(in_reg_wire_2[96])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_97
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[97]),
    .out(in_reg_wire_2[97])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_98
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[98]),
    .out(in_reg_wire_2[98])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_99
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[99]),
    .out(in_reg_wire_2[99])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_100
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[100]),
    .out(in_reg_wire_2[100])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_101
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[101]),
    .out(in_reg_wire_2[101])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_102
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[102]),
    .out(in_reg_wire_2[102])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_103
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[103]),
    .out(in_reg_wire_2[103])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_104
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[104]),
    .out(in_reg_wire_2[104])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_105
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[105]),
    .out(in_reg_wire_2[105])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_106
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[106]),
    .out(in_reg_wire_2[106])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_107
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[107]),
    .out(in_reg_wire_2[107])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_108
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[108]),
    .out(in_reg_wire_2[108])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_109
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[109]),
    .out(in_reg_wire_2[109])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_110
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[110]),
    .out(in_reg_wire_2[110])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_111
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[111]),
    .out(in_reg_wire_2[111])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_112
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[112]),
    .out(in_reg_wire_2[112])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_113
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[113]),
    .out(in_reg_wire_2[113])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_114
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[114]),
    .out(in_reg_wire_2[114])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_115
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[115]),
    .out(in_reg_wire_2[115])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_116
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[116]),
    .out(in_reg_wire_2[116])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_117
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[117]),
    .out(in_reg_wire_2[117])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_118
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[118]),
    .out(in_reg_wire_2[118])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_119
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[119]),
    .out(in_reg_wire_2[119])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_120
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[120]),
    .out(in_reg_wire_2[120])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_121
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[121]),
    .out(in_reg_wire_2[121])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_122
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[122]),
    .out(in_reg_wire_2[122])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_123
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[123]),
    .out(in_reg_wire_2[123])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_124
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[124]),
    .out(in_reg_wire_2[124])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_125
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[125]),
    .out(in_reg_wire_2[125])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_126
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[126]),
    .out(in_reg_wire_2[126])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_127
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[127]),
    .out(in_reg_wire_2[127])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_128
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[128]),
    .out(in_reg_wire_2[128])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_129
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[129]),
    .out(in_reg_wire_2[129])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_130
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[130]),
    .out(in_reg_wire_2[130])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_131
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[131]),
    .out(in_reg_wire_2[131])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_132
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[132]),
    .out(in_reg_wire_2[132])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_133
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[133]),
    .out(in_reg_wire_2[133])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_134
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[134]),
    .out(in_reg_wire_2[134])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_135
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[135]),
    .out(in_reg_wire_2[135])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_136
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[136]),
    .out(in_reg_wire_2[136])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_137
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[137]),
    .out(in_reg_wire_2[137])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_138
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[138]),
    .out(in_reg_wire_2[138])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_139
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[139]),
    .out(in_reg_wire_2[139])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_140
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[140]),
    .out(in_reg_wire_2[140])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_141
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[141]),
    .out(in_reg_wire_2[141])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_142
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[142]),
    .out(in_reg_wire_2[142])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_143
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[143]),
    .out(in_reg_wire_2[143])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_144
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[144]),
    .out(in_reg_wire_2[144])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_145
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[145]),
    .out(in_reg_wire_2[145])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_146
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[146]),
    .out(in_reg_wire_2[146])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_147
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[147]),
    .out(in_reg_wire_2[147])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_148
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[148]),
    .out(in_reg_wire_2[148])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_149
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[149]),
    .out(in_reg_wire_2[149])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_150
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[150]),
    .out(in_reg_wire_2[150])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_151
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[151]),
    .out(in_reg_wire_2[151])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_152
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[152]),
    .out(in_reg_wire_2[152])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_153
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[153]),
    .out(in_reg_wire_2[153])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_154
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[154]),
    .out(in_reg_wire_2[154])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_155
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[155]),
    .out(in_reg_wire_2[155])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_156
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[156]),
    .out(in_reg_wire_2[156])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_157
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[157]),
    .out(in_reg_wire_2[157])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_158
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[158]),
    .out(in_reg_wire_2[158])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_159
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[159]),
    .out(in_reg_wire_2[159])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_160
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[160]),
    .out(in_reg_wire_2[160])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_161
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[161]),
    .out(in_reg_wire_2[161])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_162
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[162]),
    .out(in_reg_wire_2[162])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_163
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[163]),
    .out(in_reg_wire_2[163])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_164
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[164]),
    .out(in_reg_wire_2[164])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_165
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[165]),
    .out(in_reg_wire_2[165])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_166
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[166]),
    .out(in_reg_wire_2[166])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_167
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[167]),
    .out(in_reg_wire_2[167])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_168
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[168]),
    .out(in_reg_wire_2[168])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_169
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[169]),
    .out(in_reg_wire_2[169])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_170
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[170]),
    .out(in_reg_wire_2[170])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_171
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[171]),
    .out(in_reg_wire_2[171])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_172
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[172]),
    .out(in_reg_wire_2[172])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_173
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[173]),
    .out(in_reg_wire_2[173])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_174
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[174]),
    .out(in_reg_wire_2[174])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_175
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[175]),
    .out(in_reg_wire_2[175])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_176
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[176]),
    .out(in_reg_wire_2[176])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_177
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[177]),
    .out(in_reg_wire_2[177])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_178
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[178]),
    .out(in_reg_wire_2[178])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_179
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[179]),
    .out(in_reg_wire_2[179])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_180
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[180]),
    .out(in_reg_wire_2[180])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_181
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[181]),
    .out(in_reg_wire_2[181])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_182
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[182]),
    .out(in_reg_wire_2[182])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_183
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[183]),
    .out(in_reg_wire_2[183])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_184
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[184]),
    .out(in_reg_wire_2[184])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_185
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[185]),
    .out(in_reg_wire_2[185])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_186
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[186]),
    .out(in_reg_wire_2[186])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_187
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[187]),
    .out(in_reg_wire_2[187])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_188
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[188]),
    .out(in_reg_wire_2[188])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_189
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[189]),
    .out(in_reg_wire_2[189])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_190
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[190]),
    .out(in_reg_wire_2[190])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_191
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[191]),
    .out(in_reg_wire_2[191])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_192
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[192]),
    .out(in_reg_wire_2[192])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_193
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[193]),
    .out(in_reg_wire_2[193])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_194
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[194]),
    .out(in_reg_wire_2[194])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_195
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[195]),
    .out(in_reg_wire_2[195])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_196
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[196]),
    .out(in_reg_wire_2[196])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_197
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[197]),
    .out(in_reg_wire_2[197])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_198
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[198]),
    .out(in_reg_wire_2[198])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_199
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[199]),
    .out(in_reg_wire_2[199])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_200
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[200]),
    .out(in_reg_wire_2[200])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_201
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[201]),
    .out(in_reg_wire_2[201])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_202
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[202]),
    .out(in_reg_wire_2[202])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_203
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[203]),
    .out(in_reg_wire_2[203])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_204
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[204]),
    .out(in_reg_wire_2[204])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_205
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[205]),
    .out(in_reg_wire_2[205])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_206
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[206]),
    .out(in_reg_wire_2[206])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_207
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[207]),
    .out(in_reg_wire_2[207])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_208
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[208]),
    .out(in_reg_wire_2[208])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_209
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[209]),
    .out(in_reg_wire_2[209])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_210
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[210]),
    .out(in_reg_wire_2[210])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_211
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[211]),
    .out(in_reg_wire_2[211])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_212
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[212]),
    .out(in_reg_wire_2[212])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_213
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[213]),
    .out(in_reg_wire_2[213])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_214
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[214]),
    .out(in_reg_wire_2[214])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_215
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[215]),
    .out(in_reg_wire_2[215])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_216
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[216]),
    .out(in_reg_wire_2[216])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_217
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[217]),
    .out(in_reg_wire_2[217])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_218
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[218]),
    .out(in_reg_wire_2[218])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_219
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[219]),
    .out(in_reg_wire_2[219])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_220
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[220]),
    .out(in_reg_wire_2[220])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_221
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[221]),
    .out(in_reg_wire_2[221])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_222
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[222]),
    .out(in_reg_wire_2[222])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_223
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[223]),
    .out(in_reg_wire_2[223])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_224
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[224]),
    .out(in_reg_wire_2[224])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_225
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[225]),
    .out(in_reg_wire_2[225])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_226
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[226]),
    .out(in_reg_wire_2[226])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_227
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[227]),
    .out(in_reg_wire_2[227])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_228
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[228]),
    .out(in_reg_wire_2[228])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_229
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[229]),
    .out(in_reg_wire_2[229])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_230
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[230]),
    .out(in_reg_wire_2[230])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_231
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[231]),
    .out(in_reg_wire_2[231])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_232
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[232]),
    .out(in_reg_wire_2[232])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_233
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[233]),
    .out(in_reg_wire_2[233])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_234
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[234]),
    .out(in_reg_wire_2[234])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_235
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[235]),
    .out(in_reg_wire_2[235])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_236
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[236]),
    .out(in_reg_wire_2[236])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_237
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[237]),
    .out(in_reg_wire_2[237])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_238
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[238]),
    .out(in_reg_wire_2[238])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_239
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[239]),
    .out(in_reg_wire_2[239])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_240
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[240]),
    .out(in_reg_wire_2[240])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_241
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[241]),
    .out(in_reg_wire_2[241])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_242
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[242]),
    .out(in_reg_wire_2[242])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_243
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[243]),
    .out(in_reg_wire_2[243])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_244
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[244]),
    .out(in_reg_wire_2[244])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_245
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[245]),
    .out(in_reg_wire_2[245])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_246
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[246]),
    .out(in_reg_wire_2[246])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_247
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[247]),
    .out(in_reg_wire_2[247])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_248
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[248]),
    .out(in_reg_wire_2[248])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_249
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[249]),
    .out(in_reg_wire_2[249])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_250
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[250]),
    .out(in_reg_wire_2[250])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_251
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[251]),
    .out(in_reg_wire_2[251])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_252
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[252]),
    .out(in_reg_wire_2[252])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_253
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[253]),
    .out(in_reg_wire_2[253])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_254
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[254]),
    .out(in_reg_wire_2[254])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_255
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[255]),
    .out(in_reg_wire_2[255])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_0
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[0]),
    .out(in_reg_wire_4[0])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_1
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[1]),
    .out(in_reg_wire_4[1])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_2
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[2]),
    .out(in_reg_wire_4[2])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_3
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[3]),
    .out(in_reg_wire_4[3])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_4
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[4]),
    .out(in_reg_wire_4[4])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_5
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[5]),
    .out(in_reg_wire_4[5])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_6
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[6]),
    .out(in_reg_wire_4[6])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_7
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[7]),
    .out(in_reg_wire_4[7])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_8
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[8]),
    .out(in_reg_wire_4[8])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_9
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[9]),
    .out(in_reg_wire_4[9])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_10
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[10]),
    .out(in_reg_wire_4[10])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_11
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[11]),
    .out(in_reg_wire_4[11])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_12
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[12]),
    .out(in_reg_wire_4[12])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_13
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[13]),
    .out(in_reg_wire_4[13])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_14
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[14]),
    .out(in_reg_wire_4[14])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_15
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[15]),
    .out(in_reg_wire_4[15])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_16
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[16]),
    .out(in_reg_wire_4[16])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_17
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[17]),
    .out(in_reg_wire_4[17])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_18
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[18]),
    .out(in_reg_wire_4[18])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_19
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[19]),
    .out(in_reg_wire_4[19])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_20
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[20]),
    .out(in_reg_wire_4[20])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_21
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[21]),
    .out(in_reg_wire_4[21])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_22
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[22]),
    .out(in_reg_wire_4[22])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_23
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[23]),
    .out(in_reg_wire_4[23])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_24
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[24]),
    .out(in_reg_wire_4[24])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_25
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[25]),
    .out(in_reg_wire_4[25])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_26
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[26]),
    .out(in_reg_wire_4[26])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_27
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[27]),
    .out(in_reg_wire_4[27])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_28
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[28]),
    .out(in_reg_wire_4[28])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_29
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[29]),
    .out(in_reg_wire_4[29])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_30
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[30]),
    .out(in_reg_wire_4[30])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_31
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[31]),
    .out(in_reg_wire_4[31])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_32
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[32]),
    .out(in_reg_wire_4[32])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_33
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[33]),
    .out(in_reg_wire_4[33])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_34
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[34]),
    .out(in_reg_wire_4[34])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_35
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[35]),
    .out(in_reg_wire_4[35])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_36
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[36]),
    .out(in_reg_wire_4[36])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_37
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[37]),
    .out(in_reg_wire_4[37])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_38
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[38]),
    .out(in_reg_wire_4[38])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_39
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[39]),
    .out(in_reg_wire_4[39])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_40
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[40]),
    .out(in_reg_wire_4[40])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_41
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[41]),
    .out(in_reg_wire_4[41])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_42
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[42]),
    .out(in_reg_wire_4[42])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_43
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[43]),
    .out(in_reg_wire_4[43])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_44
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[44]),
    .out(in_reg_wire_4[44])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_45
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[45]),
    .out(in_reg_wire_4[45])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_46
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[46]),
    .out(in_reg_wire_4[46])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_47
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[47]),
    .out(in_reg_wire_4[47])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_48
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[48]),
    .out(in_reg_wire_4[48])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_49
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[49]),
    .out(in_reg_wire_4[49])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_50
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[50]),
    .out(in_reg_wire_4[50])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_51
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[51]),
    .out(in_reg_wire_4[51])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_52
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[52]),
    .out(in_reg_wire_4[52])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_53
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[53]),
    .out(in_reg_wire_4[53])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_54
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[54]),
    .out(in_reg_wire_4[54])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_55
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[55]),
    .out(in_reg_wire_4[55])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_56
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[56]),
    .out(in_reg_wire_4[56])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_57
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[57]),
    .out(in_reg_wire_4[57])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_58
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[58]),
    .out(in_reg_wire_4[58])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_59
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[59]),
    .out(in_reg_wire_4[59])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_60
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[60]),
    .out(in_reg_wire_4[60])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_61
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[61]),
    .out(in_reg_wire_4[61])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_62
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[62]),
    .out(in_reg_wire_4[62])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_63
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[63]),
    .out(in_reg_wire_4[63])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_64
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[64]),
    .out(in_reg_wire_4[64])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_65
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[65]),
    .out(in_reg_wire_4[65])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_66
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[66]),
    .out(in_reg_wire_4[66])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_67
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[67]),
    .out(in_reg_wire_4[67])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_68
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[68]),
    .out(in_reg_wire_4[68])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_69
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[69]),
    .out(in_reg_wire_4[69])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_70
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[70]),
    .out(in_reg_wire_4[70])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_71
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[71]),
    .out(in_reg_wire_4[71])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_72
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[72]),
    .out(in_reg_wire_4[72])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_73
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[73]),
    .out(in_reg_wire_4[73])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_74
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[74]),
    .out(in_reg_wire_4[74])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_75
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[75]),
    .out(in_reg_wire_4[75])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_76
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[76]),
    .out(in_reg_wire_4[76])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_77
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[77]),
    .out(in_reg_wire_4[77])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_78
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[78]),
    .out(in_reg_wire_4[78])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_79
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[79]),
    .out(in_reg_wire_4[79])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_80
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[80]),
    .out(in_reg_wire_4[80])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_81
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[81]),
    .out(in_reg_wire_4[81])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_82
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[82]),
    .out(in_reg_wire_4[82])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_83
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[83]),
    .out(in_reg_wire_4[83])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_84
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[84]),
    .out(in_reg_wire_4[84])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_85
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[85]),
    .out(in_reg_wire_4[85])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_86
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[86]),
    .out(in_reg_wire_4[86])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_87
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[87]),
    .out(in_reg_wire_4[87])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_88
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[88]),
    .out(in_reg_wire_4[88])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_89
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[89]),
    .out(in_reg_wire_4[89])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_90
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[90]),
    .out(in_reg_wire_4[90])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_91
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[91]),
    .out(in_reg_wire_4[91])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_92
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[92]),
    .out(in_reg_wire_4[92])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_93
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[93]),
    .out(in_reg_wire_4[93])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_94
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[94]),
    .out(in_reg_wire_4[94])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_95
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[95]),
    .out(in_reg_wire_4[95])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_96
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[96]),
    .out(in_reg_wire_4[96])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_97
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[97]),
    .out(in_reg_wire_4[97])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_98
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[98]),
    .out(in_reg_wire_4[98])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_99
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[99]),
    .out(in_reg_wire_4[99])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_100
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[100]),
    .out(in_reg_wire_4[100])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_101
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[101]),
    .out(in_reg_wire_4[101])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_102
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[102]),
    .out(in_reg_wire_4[102])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_103
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[103]),
    .out(in_reg_wire_4[103])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_104
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[104]),
    .out(in_reg_wire_4[104])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_105
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[105]),
    .out(in_reg_wire_4[105])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_106
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[106]),
    .out(in_reg_wire_4[106])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_107
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[107]),
    .out(in_reg_wire_4[107])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_108
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[108]),
    .out(in_reg_wire_4[108])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_109
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[109]),
    .out(in_reg_wire_4[109])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_110
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[110]),
    .out(in_reg_wire_4[110])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_111
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[111]),
    .out(in_reg_wire_4[111])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_112
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[112]),
    .out(in_reg_wire_4[112])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_113
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[113]),
    .out(in_reg_wire_4[113])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_114
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[114]),
    .out(in_reg_wire_4[114])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_115
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[115]),
    .out(in_reg_wire_4[115])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_116
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[116]),
    .out(in_reg_wire_4[116])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_117
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[117]),
    .out(in_reg_wire_4[117])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_118
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[118]),
    .out(in_reg_wire_4[118])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_119
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[119]),
    .out(in_reg_wire_4[119])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_120
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[120]),
    .out(in_reg_wire_4[120])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_121
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[121]),
    .out(in_reg_wire_4[121])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_122
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[122]),
    .out(in_reg_wire_4[122])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_123
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[123]),
    .out(in_reg_wire_4[123])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_124
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[124]),
    .out(in_reg_wire_4[124])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_125
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[125]),
    .out(in_reg_wire_4[125])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_126
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[126]),
    .out(in_reg_wire_4[126])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_127
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[127]),
    .out(in_reg_wire_4[127])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_128
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[128]),
    .out(in_reg_wire_4[128])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_129
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[129]),
    .out(in_reg_wire_4[129])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_130
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[130]),
    .out(in_reg_wire_4[130])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_131
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[131]),
    .out(in_reg_wire_4[131])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_132
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[132]),
    .out(in_reg_wire_4[132])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_133
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[133]),
    .out(in_reg_wire_4[133])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_134
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[134]),
    .out(in_reg_wire_4[134])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_135
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[135]),
    .out(in_reg_wire_4[135])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_136
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[136]),
    .out(in_reg_wire_4[136])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_137
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[137]),
    .out(in_reg_wire_4[137])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_138
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[138]),
    .out(in_reg_wire_4[138])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_139
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[139]),
    .out(in_reg_wire_4[139])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_140
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[140]),
    .out(in_reg_wire_4[140])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_141
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[141]),
    .out(in_reg_wire_4[141])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_142
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[142]),
    .out(in_reg_wire_4[142])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_143
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[143]),
    .out(in_reg_wire_4[143])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_144
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[144]),
    .out(in_reg_wire_4[144])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_145
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[145]),
    .out(in_reg_wire_4[145])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_146
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[146]),
    .out(in_reg_wire_4[146])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_147
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[147]),
    .out(in_reg_wire_4[147])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_148
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[148]),
    .out(in_reg_wire_4[148])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_149
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[149]),
    .out(in_reg_wire_4[149])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_150
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[150]),
    .out(in_reg_wire_4[150])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_151
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[151]),
    .out(in_reg_wire_4[151])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_152
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[152]),
    .out(in_reg_wire_4[152])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_153
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[153]),
    .out(in_reg_wire_4[153])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_154
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[154]),
    .out(in_reg_wire_4[154])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_155
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[155]),
    .out(in_reg_wire_4[155])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_156
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[156]),
    .out(in_reg_wire_4[156])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_157
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[157]),
    .out(in_reg_wire_4[157])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_158
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[158]),
    .out(in_reg_wire_4[158])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_159
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[159]),
    .out(in_reg_wire_4[159])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_160
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[160]),
    .out(in_reg_wire_4[160])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_161
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[161]),
    .out(in_reg_wire_4[161])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_162
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[162]),
    .out(in_reg_wire_4[162])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_163
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[163]),
    .out(in_reg_wire_4[163])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_164
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[164]),
    .out(in_reg_wire_4[164])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_165
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[165]),
    .out(in_reg_wire_4[165])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_166
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[166]),
    .out(in_reg_wire_4[166])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_167
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[167]),
    .out(in_reg_wire_4[167])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_168
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[168]),
    .out(in_reg_wire_4[168])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_169
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[169]),
    .out(in_reg_wire_4[169])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_170
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[170]),
    .out(in_reg_wire_4[170])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_171
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[171]),
    .out(in_reg_wire_4[171])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_172
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[172]),
    .out(in_reg_wire_4[172])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_173
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[173]),
    .out(in_reg_wire_4[173])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_174
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[174]),
    .out(in_reg_wire_4[174])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_175
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[175]),
    .out(in_reg_wire_4[175])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_176
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[176]),
    .out(in_reg_wire_4[176])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_177
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[177]),
    .out(in_reg_wire_4[177])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_178
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[178]),
    .out(in_reg_wire_4[178])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_179
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[179]),
    .out(in_reg_wire_4[179])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_180
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[180]),
    .out(in_reg_wire_4[180])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_181
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[181]),
    .out(in_reg_wire_4[181])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_182
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[182]),
    .out(in_reg_wire_4[182])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_183
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[183]),
    .out(in_reg_wire_4[183])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_184
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[184]),
    .out(in_reg_wire_4[184])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_185
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[185]),
    .out(in_reg_wire_4[185])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_186
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[186]),
    .out(in_reg_wire_4[186])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_187
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[187]),
    .out(in_reg_wire_4[187])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_188
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[188]),
    .out(in_reg_wire_4[188])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_189
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[189]),
    .out(in_reg_wire_4[189])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_190
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[190]),
    .out(in_reg_wire_4[190])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_191
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[191]),
    .out(in_reg_wire_4[191])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_192
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[192]),
    .out(in_reg_wire_4[192])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_193
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[193]),
    .out(in_reg_wire_4[193])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_194
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[194]),
    .out(in_reg_wire_4[194])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_195
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[195]),
    .out(in_reg_wire_4[195])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_196
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[196]),
    .out(in_reg_wire_4[196])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_197
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[197]),
    .out(in_reg_wire_4[197])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_198
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[198]),
    .out(in_reg_wire_4[198])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_199
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[199]),
    .out(in_reg_wire_4[199])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_200
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[200]),
    .out(in_reg_wire_4[200])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_201
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[201]),
    .out(in_reg_wire_4[201])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_202
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[202]),
    .out(in_reg_wire_4[202])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_203
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[203]),
    .out(in_reg_wire_4[203])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_204
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[204]),
    .out(in_reg_wire_4[204])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_205
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[205]),
    .out(in_reg_wire_4[205])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_206
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[206]),
    .out(in_reg_wire_4[206])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_207
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[207]),
    .out(in_reg_wire_4[207])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_208
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[208]),
    .out(in_reg_wire_4[208])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_209
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[209]),
    .out(in_reg_wire_4[209])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_210
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[210]),
    .out(in_reg_wire_4[210])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_211
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[211]),
    .out(in_reg_wire_4[211])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_212
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[212]),
    .out(in_reg_wire_4[212])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_213
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[213]),
    .out(in_reg_wire_4[213])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_214
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[214]),
    .out(in_reg_wire_4[214])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_215
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[215]),
    .out(in_reg_wire_4[215])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_216
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[216]),
    .out(in_reg_wire_4[216])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_217
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[217]),
    .out(in_reg_wire_4[217])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_218
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[218]),
    .out(in_reg_wire_4[218])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_219
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[219]),
    .out(in_reg_wire_4[219])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_220
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[220]),
    .out(in_reg_wire_4[220])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_221
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[221]),
    .out(in_reg_wire_4[221])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_222
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[222]),
    .out(in_reg_wire_4[222])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_223
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[223]),
    .out(in_reg_wire_4[223])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_224
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[224]),
    .out(in_reg_wire_4[224])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_225
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[225]),
    .out(in_reg_wire_4[225])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_226
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[226]),
    .out(in_reg_wire_4[226])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_227
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[227]),
    .out(in_reg_wire_4[227])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_228
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[228]),
    .out(in_reg_wire_4[228])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_229
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[229]),
    .out(in_reg_wire_4[229])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_230
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[230]),
    .out(in_reg_wire_4[230])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_231
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[231]),
    .out(in_reg_wire_4[231])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_232
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[232]),
    .out(in_reg_wire_4[232])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_233
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[233]),
    .out(in_reg_wire_4[233])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_234
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[234]),
    .out(in_reg_wire_4[234])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_235
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[235]),
    .out(in_reg_wire_4[235])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_236
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[236]),
    .out(in_reg_wire_4[236])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_237
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[237]),
    .out(in_reg_wire_4[237])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_238
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[238]),
    .out(in_reg_wire_4[238])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_239
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[239]),
    .out(in_reg_wire_4[239])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_240
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[240]),
    .out(in_reg_wire_4[240])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_241
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[241]),
    .out(in_reg_wire_4[241])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_242
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[242]),
    .out(in_reg_wire_4[242])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_243
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[243]),
    .out(in_reg_wire_4[243])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_244
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[244]),
    .out(in_reg_wire_4[244])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_245
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[245]),
    .out(in_reg_wire_4[245])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_246
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[246]),
    .out(in_reg_wire_4[246])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_247
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[247]),
    .out(in_reg_wire_4[247])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_248
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[248]),
    .out(in_reg_wire_4[248])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_249
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[249]),
    .out(in_reg_wire_4[249])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_250
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[250]),
    .out(in_reg_wire_4[250])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_251
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[251]),
    .out(in_reg_wire_4[251])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_252
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[252]),
    .out(in_reg_wire_4[252])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_253
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[253]),
    .out(in_reg_wire_4[253])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_254
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[254]),
    .out(in_reg_wire_4[254])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_255
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[255]),
    .out(in_reg_wire_4[255])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_0
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[0]),
    .out(out0)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_1
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[1]),
    .out(out8)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_2
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[2]),
    .out(out16)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_3
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[3]),
    .out(out24)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_4
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[4]),
    .out(out32)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_5
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[5]),
    .out(out40)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_6
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[6]),
    .out(out48)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_7
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[7]),
    .out(out56)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_8
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[8]),
    .out(out64)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_9
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[9]),
    .out(out72)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_10
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[10]),
    .out(out80)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_11
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[11]),
    .out(out88)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_12
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[12]),
    .out(out96)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_13
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[13]),
    .out(out104)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_14
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[14]),
    .out(out112)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_15
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[15]),
    .out(out120)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_16
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[16]),
    .out(out128)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_17
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[17]),
    .out(out136)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_18
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[18]),
    .out(out144)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_19
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[19]),
    .out(out152)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_20
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[20]),
    .out(out160)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_21
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[21]),
    .out(out168)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_22
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[22]),
    .out(out176)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_23
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[23]),
    .out(out184)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_24
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[24]),
    .out(out192)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_25
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[25]),
    .out(out200)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_26
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[26]),
    .out(out208)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_27
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[27]),
    .out(out216)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_28
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[28]),
    .out(out224)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_29
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[29]),
    .out(out232)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_30
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[30]),
    .out(out240)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_31
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[31]),
    .out(out248)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_32
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[32]),
    .out(out1)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_33
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[33]),
    .out(out9)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_34
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[34]),
    .out(out17)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_35
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[35]),
    .out(out25)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_36
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[36]),
    .out(out33)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_37
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[37]),
    .out(out41)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_38
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[38]),
    .out(out49)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_39
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[39]),
    .out(out57)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_40
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[40]),
    .out(out65)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_41
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[41]),
    .out(out73)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_42
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[42]),
    .out(out81)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_43
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[43]),
    .out(out89)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_44
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[44]),
    .out(out97)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_45
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[45]),
    .out(out105)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_46
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[46]),
    .out(out113)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_47
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[47]),
    .out(out121)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_48
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[48]),
    .out(out129)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_49
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[49]),
    .out(out137)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_50
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[50]),
    .out(out145)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_51
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[51]),
    .out(out153)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_52
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[52]),
    .out(out161)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_53
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[53]),
    .out(out169)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_54
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[54]),
    .out(out177)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_55
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[55]),
    .out(out185)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_56
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[56]),
    .out(out193)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_57
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[57]),
    .out(out201)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_58
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[58]),
    .out(out209)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_59
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[59]),
    .out(out217)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_60
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[60]),
    .out(out225)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_61
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[61]),
    .out(out233)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_62
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[62]),
    .out(out241)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_63
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[63]),
    .out(out249)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_64
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[64]),
    .out(out2)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_65
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[65]),
    .out(out10)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_66
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[66]),
    .out(out18)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_67
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[67]),
    .out(out26)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_68
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[68]),
    .out(out34)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_69
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[69]),
    .out(out42)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_70
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[70]),
    .out(out50)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_71
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[71]),
    .out(out58)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_72
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[72]),
    .out(out66)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_73
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[73]),
    .out(out74)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_74
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[74]),
    .out(out82)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_75
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[75]),
    .out(out90)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_76
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[76]),
    .out(out98)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_77
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[77]),
    .out(out106)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_78
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[78]),
    .out(out114)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_79
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[79]),
    .out(out122)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_80
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[80]),
    .out(out130)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_81
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[81]),
    .out(out138)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_82
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[82]),
    .out(out146)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_83
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[83]),
    .out(out154)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_84
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[84]),
    .out(out162)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_85
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[85]),
    .out(out170)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_86
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[86]),
    .out(out178)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_87
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[87]),
    .out(out186)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_88
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[88]),
    .out(out194)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_89
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[89]),
    .out(out202)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_90
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[90]),
    .out(out210)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_91
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[91]),
    .out(out218)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_92
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[92]),
    .out(out226)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_93
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[93]),
    .out(out234)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_94
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[94]),
    .out(out242)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_95
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[95]),
    .out(out250)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_96
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[96]),
    .out(out3)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_97
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[97]),
    .out(out11)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_98
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[98]),
    .out(out19)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_99
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[99]),
    .out(out27)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_100
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[100]),
    .out(out35)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_101
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[101]),
    .out(out43)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_102
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[102]),
    .out(out51)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_103
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[103]),
    .out(out59)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_104
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[104]),
    .out(out67)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_105
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[105]),
    .out(out75)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_106
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[106]),
    .out(out83)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_107
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[107]),
    .out(out91)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_108
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[108]),
    .out(out99)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_109
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[109]),
    .out(out107)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_110
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[110]),
    .out(out115)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_111
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[111]),
    .out(out123)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_112
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[112]),
    .out(out131)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_113
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[113]),
    .out(out139)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_114
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[114]),
    .out(out147)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_115
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[115]),
    .out(out155)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_116
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[116]),
    .out(out163)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_117
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[117]),
    .out(out171)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_118
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[118]),
    .out(out179)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_119
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[119]),
    .out(out187)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_120
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[120]),
    .out(out195)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_121
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[121]),
    .out(out203)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_122
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[122]),
    .out(out211)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_123
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[123]),
    .out(out219)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_124
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[124]),
    .out(out227)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_125
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[125]),
    .out(out235)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_126
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[126]),
    .out(out243)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_127
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[127]),
    .out(out251)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_128
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[128]),
    .out(out4)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_129
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[129]),
    .out(out12)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_130
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[130]),
    .out(out20)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_131
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[131]),
    .out(out28)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_132
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[132]),
    .out(out36)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_133
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[133]),
    .out(out44)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_134
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[134]),
    .out(out52)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_135
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[135]),
    .out(out60)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_136
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[136]),
    .out(out68)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_137
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[137]),
    .out(out76)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_138
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[138]),
    .out(out84)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_139
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[139]),
    .out(out92)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_140
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[140]),
    .out(out100)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_141
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[141]),
    .out(out108)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_142
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[142]),
    .out(out116)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_143
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[143]),
    .out(out124)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_144
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[144]),
    .out(out132)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_145
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[145]),
    .out(out140)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_146
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[146]),
    .out(out148)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_147
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[147]),
    .out(out156)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_148
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[148]),
    .out(out164)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_149
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[149]),
    .out(out172)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_150
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[150]),
    .out(out180)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_151
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[151]),
    .out(out188)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_152
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[152]),
    .out(out196)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_153
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[153]),
    .out(out204)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_154
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[154]),
    .out(out212)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_155
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[155]),
    .out(out220)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_156
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[156]),
    .out(out228)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_157
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[157]),
    .out(out236)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_158
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[158]),
    .out(out244)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_159
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[159]),
    .out(out252)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_160
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[160]),
    .out(out5)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_161
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[161]),
    .out(out13)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_162
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[162]),
    .out(out21)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_163
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[163]),
    .out(out29)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_164
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[164]),
    .out(out37)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_165
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[165]),
    .out(out45)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_166
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[166]),
    .out(out53)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_167
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[167]),
    .out(out61)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_168
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[168]),
    .out(out69)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_169
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[169]),
    .out(out77)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_170
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[170]),
    .out(out85)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_171
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[171]),
    .out(out93)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_172
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[172]),
    .out(out101)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_173
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[173]),
    .out(out109)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_174
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[174]),
    .out(out117)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_175
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[175]),
    .out(out125)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_176
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[176]),
    .out(out133)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_177
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[177]),
    .out(out141)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_178
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[178]),
    .out(out149)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_179
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[179]),
    .out(out157)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_180
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[180]),
    .out(out165)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_181
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[181]),
    .out(out173)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_182
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[182]),
    .out(out181)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_183
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[183]),
    .out(out189)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_184
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[184]),
    .out(out197)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_185
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[185]),
    .out(out205)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_186
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[186]),
    .out(out213)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_187
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[187]),
    .out(out221)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_188
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[188]),
    .out(out229)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_189
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[189]),
    .out(out237)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_190
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[190]),
    .out(out245)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_191
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[191]),
    .out(out253)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_192
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[192]),
    .out(out6)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_193
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[193]),
    .out(out14)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_194
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[194]),
    .out(out22)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_195
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[195]),
    .out(out30)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_196
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[196]),
    .out(out38)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_197
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[197]),
    .out(out46)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_198
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[198]),
    .out(out54)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_199
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[199]),
    .out(out62)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_200
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[200]),
    .out(out70)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_201
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[201]),
    .out(out78)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_202
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[202]),
    .out(out86)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_203
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[203]),
    .out(out94)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_204
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[204]),
    .out(out102)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_205
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[205]),
    .out(out110)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_206
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[206]),
    .out(out118)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_207
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[207]),
    .out(out126)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_208
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[208]),
    .out(out134)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_209
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[209]),
    .out(out142)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_210
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[210]),
    .out(out150)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_211
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[211]),
    .out(out158)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_212
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[212]),
    .out(out166)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_213
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[213]),
    .out(out174)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_214
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[214]),
    .out(out182)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_215
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[215]),
    .out(out190)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_216
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[216]),
    .out(out198)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_217
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[217]),
    .out(out206)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_218
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[218]),
    .out(out214)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_219
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[219]),
    .out(out222)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_220
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[220]),
    .out(out230)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_221
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[221]),
    .out(out238)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_222
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[222]),
    .out(out246)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_223
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[223]),
    .out(out254)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_224
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[224]),
    .out(out7)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_225
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[225]),
    .out(out15)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_226
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[226]),
    .out(out23)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_227
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[227]),
    .out(out31)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_228
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[228]),
    .out(out39)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_229
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[229]),
    .out(out47)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_230
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[230]),
    .out(out55)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_231
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[231]),
    .out(out63)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_232
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[232]),
    .out(out71)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_233
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[233]),
    .out(out79)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_234
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[234]),
    .out(out87)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_235
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[235]),
    .out(out95)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_236
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[236]),
    .out(out103)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_237
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[237]),
    .out(out111)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_238
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[238]),
    .out(out119)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_239
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[239]),
    .out(out127)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_240
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[240]),
    .out(out135)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_241
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[241]),
    .out(out143)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_242
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[242]),
    .out(out151)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_243
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[243]),
    .out(out159)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_244
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[244]),
    .out(out167)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_245
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[245]),
    .out(out175)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_246
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[246]),
    .out(out183)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_247
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[247]),
    .out(out191)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_248
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[248]),
    .out(out199)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_249
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[249]),
    .out(out207)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_250
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[250]),
    .out(out215)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_251
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[251]),
    .out(out223)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_252
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[252]),
    .out(out231)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_253
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[253]),
    .out(out239)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_254
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[254]),
    .out(out247)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_255
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[255]),
    .out(out255)
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_0
  (
    .sel(conf_out[23:0]),
    .in0(in_reg_wire_0[0]),
    .in1(in_reg_wire_0[32]),
    .in2(in_reg_wire_0[64]),
    .in3(in_reg_wire_0[96]),
    .in4(in_reg_wire_0[128]),
    .in5(in_reg_wire_0[160]),
    .in6(in_reg_wire_0[192]),
    .in7(in_reg_wire_0[224]),
    .out0(in_reg_wire_1[0]),
    .out1(in_reg_wire_1[1]),
    .out2(in_reg_wire_1[2]),
    .out3(in_reg_wire_1[3]),
    .out4(in_reg_wire_1[4]),
    .out5(in_reg_wire_1[5]),
    .out6(in_reg_wire_1[6]),
    .out7(in_reg_wire_1[7])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_1
  (
    .sel(conf_out[47:24]),
    .in0(in_reg_wire_0[1]),
    .in1(in_reg_wire_0[33]),
    .in2(in_reg_wire_0[65]),
    .in3(in_reg_wire_0[97]),
    .in4(in_reg_wire_0[129]),
    .in5(in_reg_wire_0[161]),
    .in6(in_reg_wire_0[193]),
    .in7(in_reg_wire_0[225]),
    .out0(in_reg_wire_1[8]),
    .out1(in_reg_wire_1[9]),
    .out2(in_reg_wire_1[10]),
    .out3(in_reg_wire_1[11]),
    .out4(in_reg_wire_1[12]),
    .out5(in_reg_wire_1[13]),
    .out6(in_reg_wire_1[14]),
    .out7(in_reg_wire_1[15])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_2
  (
    .sel(conf_out[71:48]),
    .in0(in_reg_wire_0[2]),
    .in1(in_reg_wire_0[34]),
    .in2(in_reg_wire_0[66]),
    .in3(in_reg_wire_0[98]),
    .in4(in_reg_wire_0[130]),
    .in5(in_reg_wire_0[162]),
    .in6(in_reg_wire_0[194]),
    .in7(in_reg_wire_0[226]),
    .out0(in_reg_wire_1[16]),
    .out1(in_reg_wire_1[17]),
    .out2(in_reg_wire_1[18]),
    .out3(in_reg_wire_1[19]),
    .out4(in_reg_wire_1[20]),
    .out5(in_reg_wire_1[21]),
    .out6(in_reg_wire_1[22]),
    .out7(in_reg_wire_1[23])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_3
  (
    .sel(conf_out[95:72]),
    .in0(in_reg_wire_0[3]),
    .in1(in_reg_wire_0[35]),
    .in2(in_reg_wire_0[67]),
    .in3(in_reg_wire_0[99]),
    .in4(in_reg_wire_0[131]),
    .in5(in_reg_wire_0[163]),
    .in6(in_reg_wire_0[195]),
    .in7(in_reg_wire_0[227]),
    .out0(in_reg_wire_1[24]),
    .out1(in_reg_wire_1[25]),
    .out2(in_reg_wire_1[26]),
    .out3(in_reg_wire_1[27]),
    .out4(in_reg_wire_1[28]),
    .out5(in_reg_wire_1[29]),
    .out6(in_reg_wire_1[30]),
    .out7(in_reg_wire_1[31])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_4
  (
    .sel(conf_out[119:96]),
    .in0(in_reg_wire_0[4]),
    .in1(in_reg_wire_0[36]),
    .in2(in_reg_wire_0[68]),
    .in3(in_reg_wire_0[100]),
    .in4(in_reg_wire_0[132]),
    .in5(in_reg_wire_0[164]),
    .in6(in_reg_wire_0[196]),
    .in7(in_reg_wire_0[228]),
    .out0(in_reg_wire_1[32]),
    .out1(in_reg_wire_1[33]),
    .out2(in_reg_wire_1[34]),
    .out3(in_reg_wire_1[35]),
    .out4(in_reg_wire_1[36]),
    .out5(in_reg_wire_1[37]),
    .out6(in_reg_wire_1[38]),
    .out7(in_reg_wire_1[39])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_5
  (
    .sel(conf_out[143:120]),
    .in0(in_reg_wire_0[5]),
    .in1(in_reg_wire_0[37]),
    .in2(in_reg_wire_0[69]),
    .in3(in_reg_wire_0[101]),
    .in4(in_reg_wire_0[133]),
    .in5(in_reg_wire_0[165]),
    .in6(in_reg_wire_0[197]),
    .in7(in_reg_wire_0[229]),
    .out0(in_reg_wire_1[40]),
    .out1(in_reg_wire_1[41]),
    .out2(in_reg_wire_1[42]),
    .out3(in_reg_wire_1[43]),
    .out4(in_reg_wire_1[44]),
    .out5(in_reg_wire_1[45]),
    .out6(in_reg_wire_1[46]),
    .out7(in_reg_wire_1[47])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_6
  (
    .sel(conf_out[167:144]),
    .in0(in_reg_wire_0[6]),
    .in1(in_reg_wire_0[38]),
    .in2(in_reg_wire_0[70]),
    .in3(in_reg_wire_0[102]),
    .in4(in_reg_wire_0[134]),
    .in5(in_reg_wire_0[166]),
    .in6(in_reg_wire_0[198]),
    .in7(in_reg_wire_0[230]),
    .out0(in_reg_wire_1[48]),
    .out1(in_reg_wire_1[49]),
    .out2(in_reg_wire_1[50]),
    .out3(in_reg_wire_1[51]),
    .out4(in_reg_wire_1[52]),
    .out5(in_reg_wire_1[53]),
    .out6(in_reg_wire_1[54]),
    .out7(in_reg_wire_1[55])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_7
  (
    .sel(conf_out[191:168]),
    .in0(in_reg_wire_0[7]),
    .in1(in_reg_wire_0[39]),
    .in2(in_reg_wire_0[71]),
    .in3(in_reg_wire_0[103]),
    .in4(in_reg_wire_0[135]),
    .in5(in_reg_wire_0[167]),
    .in6(in_reg_wire_0[199]),
    .in7(in_reg_wire_0[231]),
    .out0(in_reg_wire_1[56]),
    .out1(in_reg_wire_1[57]),
    .out2(in_reg_wire_1[58]),
    .out3(in_reg_wire_1[59]),
    .out4(in_reg_wire_1[60]),
    .out5(in_reg_wire_1[61]),
    .out6(in_reg_wire_1[62]),
    .out7(in_reg_wire_1[63])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_8
  (
    .sel(conf_out[215:192]),
    .in0(in_reg_wire_0[8]),
    .in1(in_reg_wire_0[40]),
    .in2(in_reg_wire_0[72]),
    .in3(in_reg_wire_0[104]),
    .in4(in_reg_wire_0[136]),
    .in5(in_reg_wire_0[168]),
    .in6(in_reg_wire_0[200]),
    .in7(in_reg_wire_0[232]),
    .out0(in_reg_wire_1[64]),
    .out1(in_reg_wire_1[65]),
    .out2(in_reg_wire_1[66]),
    .out3(in_reg_wire_1[67]),
    .out4(in_reg_wire_1[68]),
    .out5(in_reg_wire_1[69]),
    .out6(in_reg_wire_1[70]),
    .out7(in_reg_wire_1[71])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_9
  (
    .sel(conf_out[239:216]),
    .in0(in_reg_wire_0[9]),
    .in1(in_reg_wire_0[41]),
    .in2(in_reg_wire_0[73]),
    .in3(in_reg_wire_0[105]),
    .in4(in_reg_wire_0[137]),
    .in5(in_reg_wire_0[169]),
    .in6(in_reg_wire_0[201]),
    .in7(in_reg_wire_0[233]),
    .out0(in_reg_wire_1[72]),
    .out1(in_reg_wire_1[73]),
    .out2(in_reg_wire_1[74]),
    .out3(in_reg_wire_1[75]),
    .out4(in_reg_wire_1[76]),
    .out5(in_reg_wire_1[77]),
    .out6(in_reg_wire_1[78]),
    .out7(in_reg_wire_1[79])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_10
  (
    .sel(conf_out[263:240]),
    .in0(in_reg_wire_0[10]),
    .in1(in_reg_wire_0[42]),
    .in2(in_reg_wire_0[74]),
    .in3(in_reg_wire_0[106]),
    .in4(in_reg_wire_0[138]),
    .in5(in_reg_wire_0[170]),
    .in6(in_reg_wire_0[202]),
    .in7(in_reg_wire_0[234]),
    .out0(in_reg_wire_1[80]),
    .out1(in_reg_wire_1[81]),
    .out2(in_reg_wire_1[82]),
    .out3(in_reg_wire_1[83]),
    .out4(in_reg_wire_1[84]),
    .out5(in_reg_wire_1[85]),
    .out6(in_reg_wire_1[86]),
    .out7(in_reg_wire_1[87])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_11
  (
    .sel(conf_out[287:264]),
    .in0(in_reg_wire_0[11]),
    .in1(in_reg_wire_0[43]),
    .in2(in_reg_wire_0[75]),
    .in3(in_reg_wire_0[107]),
    .in4(in_reg_wire_0[139]),
    .in5(in_reg_wire_0[171]),
    .in6(in_reg_wire_0[203]),
    .in7(in_reg_wire_0[235]),
    .out0(in_reg_wire_1[88]),
    .out1(in_reg_wire_1[89]),
    .out2(in_reg_wire_1[90]),
    .out3(in_reg_wire_1[91]),
    .out4(in_reg_wire_1[92]),
    .out5(in_reg_wire_1[93]),
    .out6(in_reg_wire_1[94]),
    .out7(in_reg_wire_1[95])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_12
  (
    .sel(conf_out[311:288]),
    .in0(in_reg_wire_0[12]),
    .in1(in_reg_wire_0[44]),
    .in2(in_reg_wire_0[76]),
    .in3(in_reg_wire_0[108]),
    .in4(in_reg_wire_0[140]),
    .in5(in_reg_wire_0[172]),
    .in6(in_reg_wire_0[204]),
    .in7(in_reg_wire_0[236]),
    .out0(in_reg_wire_1[96]),
    .out1(in_reg_wire_1[97]),
    .out2(in_reg_wire_1[98]),
    .out3(in_reg_wire_1[99]),
    .out4(in_reg_wire_1[100]),
    .out5(in_reg_wire_1[101]),
    .out6(in_reg_wire_1[102]),
    .out7(in_reg_wire_1[103])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_13
  (
    .sel(conf_out[335:312]),
    .in0(in_reg_wire_0[13]),
    .in1(in_reg_wire_0[45]),
    .in2(in_reg_wire_0[77]),
    .in3(in_reg_wire_0[109]),
    .in4(in_reg_wire_0[141]),
    .in5(in_reg_wire_0[173]),
    .in6(in_reg_wire_0[205]),
    .in7(in_reg_wire_0[237]),
    .out0(in_reg_wire_1[104]),
    .out1(in_reg_wire_1[105]),
    .out2(in_reg_wire_1[106]),
    .out3(in_reg_wire_1[107]),
    .out4(in_reg_wire_1[108]),
    .out5(in_reg_wire_1[109]),
    .out6(in_reg_wire_1[110]),
    .out7(in_reg_wire_1[111])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_14
  (
    .sel(conf_out[359:336]),
    .in0(in_reg_wire_0[14]),
    .in1(in_reg_wire_0[46]),
    .in2(in_reg_wire_0[78]),
    .in3(in_reg_wire_0[110]),
    .in4(in_reg_wire_0[142]),
    .in5(in_reg_wire_0[174]),
    .in6(in_reg_wire_0[206]),
    .in7(in_reg_wire_0[238]),
    .out0(in_reg_wire_1[112]),
    .out1(in_reg_wire_1[113]),
    .out2(in_reg_wire_1[114]),
    .out3(in_reg_wire_1[115]),
    .out4(in_reg_wire_1[116]),
    .out5(in_reg_wire_1[117]),
    .out6(in_reg_wire_1[118]),
    .out7(in_reg_wire_1[119])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_15
  (
    .sel(conf_out[383:360]),
    .in0(in_reg_wire_0[15]),
    .in1(in_reg_wire_0[47]),
    .in2(in_reg_wire_0[79]),
    .in3(in_reg_wire_0[111]),
    .in4(in_reg_wire_0[143]),
    .in5(in_reg_wire_0[175]),
    .in6(in_reg_wire_0[207]),
    .in7(in_reg_wire_0[239]),
    .out0(in_reg_wire_1[120]),
    .out1(in_reg_wire_1[121]),
    .out2(in_reg_wire_1[122]),
    .out3(in_reg_wire_1[123]),
    .out4(in_reg_wire_1[124]),
    .out5(in_reg_wire_1[125]),
    .out6(in_reg_wire_1[126]),
    .out7(in_reg_wire_1[127])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_16
  (
    .sel(conf_out[407:384]),
    .in0(in_reg_wire_0[16]),
    .in1(in_reg_wire_0[48]),
    .in2(in_reg_wire_0[80]),
    .in3(in_reg_wire_0[112]),
    .in4(in_reg_wire_0[144]),
    .in5(in_reg_wire_0[176]),
    .in6(in_reg_wire_0[208]),
    .in7(in_reg_wire_0[240]),
    .out0(in_reg_wire_1[128]),
    .out1(in_reg_wire_1[129]),
    .out2(in_reg_wire_1[130]),
    .out3(in_reg_wire_1[131]),
    .out4(in_reg_wire_1[132]),
    .out5(in_reg_wire_1[133]),
    .out6(in_reg_wire_1[134]),
    .out7(in_reg_wire_1[135])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_17
  (
    .sel(conf_out[431:408]),
    .in0(in_reg_wire_0[17]),
    .in1(in_reg_wire_0[49]),
    .in2(in_reg_wire_0[81]),
    .in3(in_reg_wire_0[113]),
    .in4(in_reg_wire_0[145]),
    .in5(in_reg_wire_0[177]),
    .in6(in_reg_wire_0[209]),
    .in7(in_reg_wire_0[241]),
    .out0(in_reg_wire_1[136]),
    .out1(in_reg_wire_1[137]),
    .out2(in_reg_wire_1[138]),
    .out3(in_reg_wire_1[139]),
    .out4(in_reg_wire_1[140]),
    .out5(in_reg_wire_1[141]),
    .out6(in_reg_wire_1[142]),
    .out7(in_reg_wire_1[143])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_18
  (
    .sel(conf_out[455:432]),
    .in0(in_reg_wire_0[18]),
    .in1(in_reg_wire_0[50]),
    .in2(in_reg_wire_0[82]),
    .in3(in_reg_wire_0[114]),
    .in4(in_reg_wire_0[146]),
    .in5(in_reg_wire_0[178]),
    .in6(in_reg_wire_0[210]),
    .in7(in_reg_wire_0[242]),
    .out0(in_reg_wire_1[144]),
    .out1(in_reg_wire_1[145]),
    .out2(in_reg_wire_1[146]),
    .out3(in_reg_wire_1[147]),
    .out4(in_reg_wire_1[148]),
    .out5(in_reg_wire_1[149]),
    .out6(in_reg_wire_1[150]),
    .out7(in_reg_wire_1[151])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_19
  (
    .sel(conf_out[479:456]),
    .in0(in_reg_wire_0[19]),
    .in1(in_reg_wire_0[51]),
    .in2(in_reg_wire_0[83]),
    .in3(in_reg_wire_0[115]),
    .in4(in_reg_wire_0[147]),
    .in5(in_reg_wire_0[179]),
    .in6(in_reg_wire_0[211]),
    .in7(in_reg_wire_0[243]),
    .out0(in_reg_wire_1[152]),
    .out1(in_reg_wire_1[153]),
    .out2(in_reg_wire_1[154]),
    .out3(in_reg_wire_1[155]),
    .out4(in_reg_wire_1[156]),
    .out5(in_reg_wire_1[157]),
    .out6(in_reg_wire_1[158]),
    .out7(in_reg_wire_1[159])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_20
  (
    .sel(conf_out[503:480]),
    .in0(in_reg_wire_0[20]),
    .in1(in_reg_wire_0[52]),
    .in2(in_reg_wire_0[84]),
    .in3(in_reg_wire_0[116]),
    .in4(in_reg_wire_0[148]),
    .in5(in_reg_wire_0[180]),
    .in6(in_reg_wire_0[212]),
    .in7(in_reg_wire_0[244]),
    .out0(in_reg_wire_1[160]),
    .out1(in_reg_wire_1[161]),
    .out2(in_reg_wire_1[162]),
    .out3(in_reg_wire_1[163]),
    .out4(in_reg_wire_1[164]),
    .out5(in_reg_wire_1[165]),
    .out6(in_reg_wire_1[166]),
    .out7(in_reg_wire_1[167])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_21
  (
    .sel(conf_out[527:504]),
    .in0(in_reg_wire_0[21]),
    .in1(in_reg_wire_0[53]),
    .in2(in_reg_wire_0[85]),
    .in3(in_reg_wire_0[117]),
    .in4(in_reg_wire_0[149]),
    .in5(in_reg_wire_0[181]),
    .in6(in_reg_wire_0[213]),
    .in7(in_reg_wire_0[245]),
    .out0(in_reg_wire_1[168]),
    .out1(in_reg_wire_1[169]),
    .out2(in_reg_wire_1[170]),
    .out3(in_reg_wire_1[171]),
    .out4(in_reg_wire_1[172]),
    .out5(in_reg_wire_1[173]),
    .out6(in_reg_wire_1[174]),
    .out7(in_reg_wire_1[175])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_22
  (
    .sel(conf_out[551:528]),
    .in0(in_reg_wire_0[22]),
    .in1(in_reg_wire_0[54]),
    .in2(in_reg_wire_0[86]),
    .in3(in_reg_wire_0[118]),
    .in4(in_reg_wire_0[150]),
    .in5(in_reg_wire_0[182]),
    .in6(in_reg_wire_0[214]),
    .in7(in_reg_wire_0[246]),
    .out0(in_reg_wire_1[176]),
    .out1(in_reg_wire_1[177]),
    .out2(in_reg_wire_1[178]),
    .out3(in_reg_wire_1[179]),
    .out4(in_reg_wire_1[180]),
    .out5(in_reg_wire_1[181]),
    .out6(in_reg_wire_1[182]),
    .out7(in_reg_wire_1[183])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_23
  (
    .sel(conf_out[575:552]),
    .in0(in_reg_wire_0[23]),
    .in1(in_reg_wire_0[55]),
    .in2(in_reg_wire_0[87]),
    .in3(in_reg_wire_0[119]),
    .in4(in_reg_wire_0[151]),
    .in5(in_reg_wire_0[183]),
    .in6(in_reg_wire_0[215]),
    .in7(in_reg_wire_0[247]),
    .out0(in_reg_wire_1[184]),
    .out1(in_reg_wire_1[185]),
    .out2(in_reg_wire_1[186]),
    .out3(in_reg_wire_1[187]),
    .out4(in_reg_wire_1[188]),
    .out5(in_reg_wire_1[189]),
    .out6(in_reg_wire_1[190]),
    .out7(in_reg_wire_1[191])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_24
  (
    .sel(conf_out[599:576]),
    .in0(in_reg_wire_0[24]),
    .in1(in_reg_wire_0[56]),
    .in2(in_reg_wire_0[88]),
    .in3(in_reg_wire_0[120]),
    .in4(in_reg_wire_0[152]),
    .in5(in_reg_wire_0[184]),
    .in6(in_reg_wire_0[216]),
    .in7(in_reg_wire_0[248]),
    .out0(in_reg_wire_1[192]),
    .out1(in_reg_wire_1[193]),
    .out2(in_reg_wire_1[194]),
    .out3(in_reg_wire_1[195]),
    .out4(in_reg_wire_1[196]),
    .out5(in_reg_wire_1[197]),
    .out6(in_reg_wire_1[198]),
    .out7(in_reg_wire_1[199])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_25
  (
    .sel(conf_out[623:600]),
    .in0(in_reg_wire_0[25]),
    .in1(in_reg_wire_0[57]),
    .in2(in_reg_wire_0[89]),
    .in3(in_reg_wire_0[121]),
    .in4(in_reg_wire_0[153]),
    .in5(in_reg_wire_0[185]),
    .in6(in_reg_wire_0[217]),
    .in7(in_reg_wire_0[249]),
    .out0(in_reg_wire_1[200]),
    .out1(in_reg_wire_1[201]),
    .out2(in_reg_wire_1[202]),
    .out3(in_reg_wire_1[203]),
    .out4(in_reg_wire_1[204]),
    .out5(in_reg_wire_1[205]),
    .out6(in_reg_wire_1[206]),
    .out7(in_reg_wire_1[207])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_26
  (
    .sel(conf_out[647:624]),
    .in0(in_reg_wire_0[26]),
    .in1(in_reg_wire_0[58]),
    .in2(in_reg_wire_0[90]),
    .in3(in_reg_wire_0[122]),
    .in4(in_reg_wire_0[154]),
    .in5(in_reg_wire_0[186]),
    .in6(in_reg_wire_0[218]),
    .in7(in_reg_wire_0[250]),
    .out0(in_reg_wire_1[208]),
    .out1(in_reg_wire_1[209]),
    .out2(in_reg_wire_1[210]),
    .out3(in_reg_wire_1[211]),
    .out4(in_reg_wire_1[212]),
    .out5(in_reg_wire_1[213]),
    .out6(in_reg_wire_1[214]),
    .out7(in_reg_wire_1[215])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_27
  (
    .sel(conf_out[671:648]),
    .in0(in_reg_wire_0[27]),
    .in1(in_reg_wire_0[59]),
    .in2(in_reg_wire_0[91]),
    .in3(in_reg_wire_0[123]),
    .in4(in_reg_wire_0[155]),
    .in5(in_reg_wire_0[187]),
    .in6(in_reg_wire_0[219]),
    .in7(in_reg_wire_0[251]),
    .out0(in_reg_wire_1[216]),
    .out1(in_reg_wire_1[217]),
    .out2(in_reg_wire_1[218]),
    .out3(in_reg_wire_1[219]),
    .out4(in_reg_wire_1[220]),
    .out5(in_reg_wire_1[221]),
    .out6(in_reg_wire_1[222]),
    .out7(in_reg_wire_1[223])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_28
  (
    .sel(conf_out[695:672]),
    .in0(in_reg_wire_0[28]),
    .in1(in_reg_wire_0[60]),
    .in2(in_reg_wire_0[92]),
    .in3(in_reg_wire_0[124]),
    .in4(in_reg_wire_0[156]),
    .in5(in_reg_wire_0[188]),
    .in6(in_reg_wire_0[220]),
    .in7(in_reg_wire_0[252]),
    .out0(in_reg_wire_1[224]),
    .out1(in_reg_wire_1[225]),
    .out2(in_reg_wire_1[226]),
    .out3(in_reg_wire_1[227]),
    .out4(in_reg_wire_1[228]),
    .out5(in_reg_wire_1[229]),
    .out6(in_reg_wire_1[230]),
    .out7(in_reg_wire_1[231])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_29
  (
    .sel(conf_out[719:696]),
    .in0(in_reg_wire_0[29]),
    .in1(in_reg_wire_0[61]),
    .in2(in_reg_wire_0[93]),
    .in3(in_reg_wire_0[125]),
    .in4(in_reg_wire_0[157]),
    .in5(in_reg_wire_0[189]),
    .in6(in_reg_wire_0[221]),
    .in7(in_reg_wire_0[253]),
    .out0(in_reg_wire_1[232]),
    .out1(in_reg_wire_1[233]),
    .out2(in_reg_wire_1[234]),
    .out3(in_reg_wire_1[235]),
    .out4(in_reg_wire_1[236]),
    .out5(in_reg_wire_1[237]),
    .out6(in_reg_wire_1[238]),
    .out7(in_reg_wire_1[239])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_30
  (
    .sel(conf_out[743:720]),
    .in0(in_reg_wire_0[30]),
    .in1(in_reg_wire_0[62]),
    .in2(in_reg_wire_0[94]),
    .in3(in_reg_wire_0[126]),
    .in4(in_reg_wire_0[158]),
    .in5(in_reg_wire_0[190]),
    .in6(in_reg_wire_0[222]),
    .in7(in_reg_wire_0[254]),
    .out0(in_reg_wire_1[240]),
    .out1(in_reg_wire_1[241]),
    .out2(in_reg_wire_1[242]),
    .out3(in_reg_wire_1[243]),
    .out4(in_reg_wire_1[244]),
    .out5(in_reg_wire_1[245]),
    .out6(in_reg_wire_1[246]),
    .out7(in_reg_wire_1[247])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_31
  (
    .sel(conf_out[767:744]),
    .in0(in_reg_wire_0[31]),
    .in1(in_reg_wire_0[63]),
    .in2(in_reg_wire_0[95]),
    .in3(in_reg_wire_0[127]),
    .in4(in_reg_wire_0[159]),
    .in5(in_reg_wire_0[191]),
    .in6(in_reg_wire_0[223]),
    .in7(in_reg_wire_0[255]),
    .out0(in_reg_wire_1[248]),
    .out1(in_reg_wire_1[249]),
    .out2(in_reg_wire_1[250]),
    .out3(in_reg_wire_1[251]),
    .out4(in_reg_wire_1[252]),
    .out5(in_reg_wire_1[253]),
    .out6(in_reg_wire_1[254]),
    .out7(in_reg_wire_1[255])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_0
  (
    .sel(conf_out[791:768]),
    .in0(in_reg_wire_2[0]),
    .in1(in_reg_wire_2[32]),
    .in2(in_reg_wire_2[64]),
    .in3(in_reg_wire_2[96]),
    .in4(in_reg_wire_2[128]),
    .in5(in_reg_wire_2[160]),
    .in6(in_reg_wire_2[192]),
    .in7(in_reg_wire_2[224]),
    .out0(in_reg_wire_3[0]),
    .out1(in_reg_wire_3[1]),
    .out2(in_reg_wire_3[2]),
    .out3(in_reg_wire_3[3]),
    .out4(in_reg_wire_3[4]),
    .out5(in_reg_wire_3[5]),
    .out6(in_reg_wire_3[6]),
    .out7(in_reg_wire_3[7])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_1
  (
    .sel(conf_out[815:792]),
    .in0(in_reg_wire_2[1]),
    .in1(in_reg_wire_2[33]),
    .in2(in_reg_wire_2[65]),
    .in3(in_reg_wire_2[97]),
    .in4(in_reg_wire_2[129]),
    .in5(in_reg_wire_2[161]),
    .in6(in_reg_wire_2[193]),
    .in7(in_reg_wire_2[225]),
    .out0(in_reg_wire_3[8]),
    .out1(in_reg_wire_3[9]),
    .out2(in_reg_wire_3[10]),
    .out3(in_reg_wire_3[11]),
    .out4(in_reg_wire_3[12]),
    .out5(in_reg_wire_3[13]),
    .out6(in_reg_wire_3[14]),
    .out7(in_reg_wire_3[15])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_2
  (
    .sel(conf_out[839:816]),
    .in0(in_reg_wire_2[2]),
    .in1(in_reg_wire_2[34]),
    .in2(in_reg_wire_2[66]),
    .in3(in_reg_wire_2[98]),
    .in4(in_reg_wire_2[130]),
    .in5(in_reg_wire_2[162]),
    .in6(in_reg_wire_2[194]),
    .in7(in_reg_wire_2[226]),
    .out0(in_reg_wire_3[16]),
    .out1(in_reg_wire_3[17]),
    .out2(in_reg_wire_3[18]),
    .out3(in_reg_wire_3[19]),
    .out4(in_reg_wire_3[20]),
    .out5(in_reg_wire_3[21]),
    .out6(in_reg_wire_3[22]),
    .out7(in_reg_wire_3[23])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_3
  (
    .sel(conf_out[863:840]),
    .in0(in_reg_wire_2[3]),
    .in1(in_reg_wire_2[35]),
    .in2(in_reg_wire_2[67]),
    .in3(in_reg_wire_2[99]),
    .in4(in_reg_wire_2[131]),
    .in5(in_reg_wire_2[163]),
    .in6(in_reg_wire_2[195]),
    .in7(in_reg_wire_2[227]),
    .out0(in_reg_wire_3[24]),
    .out1(in_reg_wire_3[25]),
    .out2(in_reg_wire_3[26]),
    .out3(in_reg_wire_3[27]),
    .out4(in_reg_wire_3[28]),
    .out5(in_reg_wire_3[29]),
    .out6(in_reg_wire_3[30]),
    .out7(in_reg_wire_3[31])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_4
  (
    .sel(conf_out[887:864]),
    .in0(in_reg_wire_2[4]),
    .in1(in_reg_wire_2[36]),
    .in2(in_reg_wire_2[68]),
    .in3(in_reg_wire_2[100]),
    .in4(in_reg_wire_2[132]),
    .in5(in_reg_wire_2[164]),
    .in6(in_reg_wire_2[196]),
    .in7(in_reg_wire_2[228]),
    .out0(in_reg_wire_3[32]),
    .out1(in_reg_wire_3[33]),
    .out2(in_reg_wire_3[34]),
    .out3(in_reg_wire_3[35]),
    .out4(in_reg_wire_3[36]),
    .out5(in_reg_wire_3[37]),
    .out6(in_reg_wire_3[38]),
    .out7(in_reg_wire_3[39])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_5
  (
    .sel(conf_out[911:888]),
    .in0(in_reg_wire_2[5]),
    .in1(in_reg_wire_2[37]),
    .in2(in_reg_wire_2[69]),
    .in3(in_reg_wire_2[101]),
    .in4(in_reg_wire_2[133]),
    .in5(in_reg_wire_2[165]),
    .in6(in_reg_wire_2[197]),
    .in7(in_reg_wire_2[229]),
    .out0(in_reg_wire_3[40]),
    .out1(in_reg_wire_3[41]),
    .out2(in_reg_wire_3[42]),
    .out3(in_reg_wire_3[43]),
    .out4(in_reg_wire_3[44]),
    .out5(in_reg_wire_3[45]),
    .out6(in_reg_wire_3[46]),
    .out7(in_reg_wire_3[47])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_6
  (
    .sel(conf_out[935:912]),
    .in0(in_reg_wire_2[6]),
    .in1(in_reg_wire_2[38]),
    .in2(in_reg_wire_2[70]),
    .in3(in_reg_wire_2[102]),
    .in4(in_reg_wire_2[134]),
    .in5(in_reg_wire_2[166]),
    .in6(in_reg_wire_2[198]),
    .in7(in_reg_wire_2[230]),
    .out0(in_reg_wire_3[48]),
    .out1(in_reg_wire_3[49]),
    .out2(in_reg_wire_3[50]),
    .out3(in_reg_wire_3[51]),
    .out4(in_reg_wire_3[52]),
    .out5(in_reg_wire_3[53]),
    .out6(in_reg_wire_3[54]),
    .out7(in_reg_wire_3[55])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_7
  (
    .sel(conf_out[959:936]),
    .in0(in_reg_wire_2[7]),
    .in1(in_reg_wire_2[39]),
    .in2(in_reg_wire_2[71]),
    .in3(in_reg_wire_2[103]),
    .in4(in_reg_wire_2[135]),
    .in5(in_reg_wire_2[167]),
    .in6(in_reg_wire_2[199]),
    .in7(in_reg_wire_2[231]),
    .out0(in_reg_wire_3[56]),
    .out1(in_reg_wire_3[57]),
    .out2(in_reg_wire_3[58]),
    .out3(in_reg_wire_3[59]),
    .out4(in_reg_wire_3[60]),
    .out5(in_reg_wire_3[61]),
    .out6(in_reg_wire_3[62]),
    .out7(in_reg_wire_3[63])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_8
  (
    .sel(conf_out[983:960]),
    .in0(in_reg_wire_2[8]),
    .in1(in_reg_wire_2[40]),
    .in2(in_reg_wire_2[72]),
    .in3(in_reg_wire_2[104]),
    .in4(in_reg_wire_2[136]),
    .in5(in_reg_wire_2[168]),
    .in6(in_reg_wire_2[200]),
    .in7(in_reg_wire_2[232]),
    .out0(in_reg_wire_3[64]),
    .out1(in_reg_wire_3[65]),
    .out2(in_reg_wire_3[66]),
    .out3(in_reg_wire_3[67]),
    .out4(in_reg_wire_3[68]),
    .out5(in_reg_wire_3[69]),
    .out6(in_reg_wire_3[70]),
    .out7(in_reg_wire_3[71])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_9
  (
    .sel(conf_out[1007:984]),
    .in0(in_reg_wire_2[9]),
    .in1(in_reg_wire_2[41]),
    .in2(in_reg_wire_2[73]),
    .in3(in_reg_wire_2[105]),
    .in4(in_reg_wire_2[137]),
    .in5(in_reg_wire_2[169]),
    .in6(in_reg_wire_2[201]),
    .in7(in_reg_wire_2[233]),
    .out0(in_reg_wire_3[72]),
    .out1(in_reg_wire_3[73]),
    .out2(in_reg_wire_3[74]),
    .out3(in_reg_wire_3[75]),
    .out4(in_reg_wire_3[76]),
    .out5(in_reg_wire_3[77]),
    .out6(in_reg_wire_3[78]),
    .out7(in_reg_wire_3[79])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_10
  (
    .sel(conf_out[1031:1008]),
    .in0(in_reg_wire_2[10]),
    .in1(in_reg_wire_2[42]),
    .in2(in_reg_wire_2[74]),
    .in3(in_reg_wire_2[106]),
    .in4(in_reg_wire_2[138]),
    .in5(in_reg_wire_2[170]),
    .in6(in_reg_wire_2[202]),
    .in7(in_reg_wire_2[234]),
    .out0(in_reg_wire_3[80]),
    .out1(in_reg_wire_3[81]),
    .out2(in_reg_wire_3[82]),
    .out3(in_reg_wire_3[83]),
    .out4(in_reg_wire_3[84]),
    .out5(in_reg_wire_3[85]),
    .out6(in_reg_wire_3[86]),
    .out7(in_reg_wire_3[87])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_11
  (
    .sel(conf_out[1055:1032]),
    .in0(in_reg_wire_2[11]),
    .in1(in_reg_wire_2[43]),
    .in2(in_reg_wire_2[75]),
    .in3(in_reg_wire_2[107]),
    .in4(in_reg_wire_2[139]),
    .in5(in_reg_wire_2[171]),
    .in6(in_reg_wire_2[203]),
    .in7(in_reg_wire_2[235]),
    .out0(in_reg_wire_3[88]),
    .out1(in_reg_wire_3[89]),
    .out2(in_reg_wire_3[90]),
    .out3(in_reg_wire_3[91]),
    .out4(in_reg_wire_3[92]),
    .out5(in_reg_wire_3[93]),
    .out6(in_reg_wire_3[94]),
    .out7(in_reg_wire_3[95])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_12
  (
    .sel(conf_out[1079:1056]),
    .in0(in_reg_wire_2[12]),
    .in1(in_reg_wire_2[44]),
    .in2(in_reg_wire_2[76]),
    .in3(in_reg_wire_2[108]),
    .in4(in_reg_wire_2[140]),
    .in5(in_reg_wire_2[172]),
    .in6(in_reg_wire_2[204]),
    .in7(in_reg_wire_2[236]),
    .out0(in_reg_wire_3[96]),
    .out1(in_reg_wire_3[97]),
    .out2(in_reg_wire_3[98]),
    .out3(in_reg_wire_3[99]),
    .out4(in_reg_wire_3[100]),
    .out5(in_reg_wire_3[101]),
    .out6(in_reg_wire_3[102]),
    .out7(in_reg_wire_3[103])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_13
  (
    .sel(conf_out[1103:1080]),
    .in0(in_reg_wire_2[13]),
    .in1(in_reg_wire_2[45]),
    .in2(in_reg_wire_2[77]),
    .in3(in_reg_wire_2[109]),
    .in4(in_reg_wire_2[141]),
    .in5(in_reg_wire_2[173]),
    .in6(in_reg_wire_2[205]),
    .in7(in_reg_wire_2[237]),
    .out0(in_reg_wire_3[104]),
    .out1(in_reg_wire_3[105]),
    .out2(in_reg_wire_3[106]),
    .out3(in_reg_wire_3[107]),
    .out4(in_reg_wire_3[108]),
    .out5(in_reg_wire_3[109]),
    .out6(in_reg_wire_3[110]),
    .out7(in_reg_wire_3[111])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_14
  (
    .sel(conf_out[1127:1104]),
    .in0(in_reg_wire_2[14]),
    .in1(in_reg_wire_2[46]),
    .in2(in_reg_wire_2[78]),
    .in3(in_reg_wire_2[110]),
    .in4(in_reg_wire_2[142]),
    .in5(in_reg_wire_2[174]),
    .in6(in_reg_wire_2[206]),
    .in7(in_reg_wire_2[238]),
    .out0(in_reg_wire_3[112]),
    .out1(in_reg_wire_3[113]),
    .out2(in_reg_wire_3[114]),
    .out3(in_reg_wire_3[115]),
    .out4(in_reg_wire_3[116]),
    .out5(in_reg_wire_3[117]),
    .out6(in_reg_wire_3[118]),
    .out7(in_reg_wire_3[119])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_15
  (
    .sel(conf_out[1151:1128]),
    .in0(in_reg_wire_2[15]),
    .in1(in_reg_wire_2[47]),
    .in2(in_reg_wire_2[79]),
    .in3(in_reg_wire_2[111]),
    .in4(in_reg_wire_2[143]),
    .in5(in_reg_wire_2[175]),
    .in6(in_reg_wire_2[207]),
    .in7(in_reg_wire_2[239]),
    .out0(in_reg_wire_3[120]),
    .out1(in_reg_wire_3[121]),
    .out2(in_reg_wire_3[122]),
    .out3(in_reg_wire_3[123]),
    .out4(in_reg_wire_3[124]),
    .out5(in_reg_wire_3[125]),
    .out6(in_reg_wire_3[126]),
    .out7(in_reg_wire_3[127])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_16
  (
    .sel(conf_out[1175:1152]),
    .in0(in_reg_wire_2[16]),
    .in1(in_reg_wire_2[48]),
    .in2(in_reg_wire_2[80]),
    .in3(in_reg_wire_2[112]),
    .in4(in_reg_wire_2[144]),
    .in5(in_reg_wire_2[176]),
    .in6(in_reg_wire_2[208]),
    .in7(in_reg_wire_2[240]),
    .out0(in_reg_wire_3[128]),
    .out1(in_reg_wire_3[129]),
    .out2(in_reg_wire_3[130]),
    .out3(in_reg_wire_3[131]),
    .out4(in_reg_wire_3[132]),
    .out5(in_reg_wire_3[133]),
    .out6(in_reg_wire_3[134]),
    .out7(in_reg_wire_3[135])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_17
  (
    .sel(conf_out[1199:1176]),
    .in0(in_reg_wire_2[17]),
    .in1(in_reg_wire_2[49]),
    .in2(in_reg_wire_2[81]),
    .in3(in_reg_wire_2[113]),
    .in4(in_reg_wire_2[145]),
    .in5(in_reg_wire_2[177]),
    .in6(in_reg_wire_2[209]),
    .in7(in_reg_wire_2[241]),
    .out0(in_reg_wire_3[136]),
    .out1(in_reg_wire_3[137]),
    .out2(in_reg_wire_3[138]),
    .out3(in_reg_wire_3[139]),
    .out4(in_reg_wire_3[140]),
    .out5(in_reg_wire_3[141]),
    .out6(in_reg_wire_3[142]),
    .out7(in_reg_wire_3[143])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_18
  (
    .sel(conf_out[1223:1200]),
    .in0(in_reg_wire_2[18]),
    .in1(in_reg_wire_2[50]),
    .in2(in_reg_wire_2[82]),
    .in3(in_reg_wire_2[114]),
    .in4(in_reg_wire_2[146]),
    .in5(in_reg_wire_2[178]),
    .in6(in_reg_wire_2[210]),
    .in7(in_reg_wire_2[242]),
    .out0(in_reg_wire_3[144]),
    .out1(in_reg_wire_3[145]),
    .out2(in_reg_wire_3[146]),
    .out3(in_reg_wire_3[147]),
    .out4(in_reg_wire_3[148]),
    .out5(in_reg_wire_3[149]),
    .out6(in_reg_wire_3[150]),
    .out7(in_reg_wire_3[151])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_19
  (
    .sel(conf_out[1247:1224]),
    .in0(in_reg_wire_2[19]),
    .in1(in_reg_wire_2[51]),
    .in2(in_reg_wire_2[83]),
    .in3(in_reg_wire_2[115]),
    .in4(in_reg_wire_2[147]),
    .in5(in_reg_wire_2[179]),
    .in6(in_reg_wire_2[211]),
    .in7(in_reg_wire_2[243]),
    .out0(in_reg_wire_3[152]),
    .out1(in_reg_wire_3[153]),
    .out2(in_reg_wire_3[154]),
    .out3(in_reg_wire_3[155]),
    .out4(in_reg_wire_3[156]),
    .out5(in_reg_wire_3[157]),
    .out6(in_reg_wire_3[158]),
    .out7(in_reg_wire_3[159])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_20
  (
    .sel(conf_out[1271:1248]),
    .in0(in_reg_wire_2[20]),
    .in1(in_reg_wire_2[52]),
    .in2(in_reg_wire_2[84]),
    .in3(in_reg_wire_2[116]),
    .in4(in_reg_wire_2[148]),
    .in5(in_reg_wire_2[180]),
    .in6(in_reg_wire_2[212]),
    .in7(in_reg_wire_2[244]),
    .out0(in_reg_wire_3[160]),
    .out1(in_reg_wire_3[161]),
    .out2(in_reg_wire_3[162]),
    .out3(in_reg_wire_3[163]),
    .out4(in_reg_wire_3[164]),
    .out5(in_reg_wire_3[165]),
    .out6(in_reg_wire_3[166]),
    .out7(in_reg_wire_3[167])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_21
  (
    .sel(conf_out[1295:1272]),
    .in0(in_reg_wire_2[21]),
    .in1(in_reg_wire_2[53]),
    .in2(in_reg_wire_2[85]),
    .in3(in_reg_wire_2[117]),
    .in4(in_reg_wire_2[149]),
    .in5(in_reg_wire_2[181]),
    .in6(in_reg_wire_2[213]),
    .in7(in_reg_wire_2[245]),
    .out0(in_reg_wire_3[168]),
    .out1(in_reg_wire_3[169]),
    .out2(in_reg_wire_3[170]),
    .out3(in_reg_wire_3[171]),
    .out4(in_reg_wire_3[172]),
    .out5(in_reg_wire_3[173]),
    .out6(in_reg_wire_3[174]),
    .out7(in_reg_wire_3[175])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_22
  (
    .sel(conf_out[1319:1296]),
    .in0(in_reg_wire_2[22]),
    .in1(in_reg_wire_2[54]),
    .in2(in_reg_wire_2[86]),
    .in3(in_reg_wire_2[118]),
    .in4(in_reg_wire_2[150]),
    .in5(in_reg_wire_2[182]),
    .in6(in_reg_wire_2[214]),
    .in7(in_reg_wire_2[246]),
    .out0(in_reg_wire_3[176]),
    .out1(in_reg_wire_3[177]),
    .out2(in_reg_wire_3[178]),
    .out3(in_reg_wire_3[179]),
    .out4(in_reg_wire_3[180]),
    .out5(in_reg_wire_3[181]),
    .out6(in_reg_wire_3[182]),
    .out7(in_reg_wire_3[183])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_23
  (
    .sel(conf_out[1343:1320]),
    .in0(in_reg_wire_2[23]),
    .in1(in_reg_wire_2[55]),
    .in2(in_reg_wire_2[87]),
    .in3(in_reg_wire_2[119]),
    .in4(in_reg_wire_2[151]),
    .in5(in_reg_wire_2[183]),
    .in6(in_reg_wire_2[215]),
    .in7(in_reg_wire_2[247]),
    .out0(in_reg_wire_3[184]),
    .out1(in_reg_wire_3[185]),
    .out2(in_reg_wire_3[186]),
    .out3(in_reg_wire_3[187]),
    .out4(in_reg_wire_3[188]),
    .out5(in_reg_wire_3[189]),
    .out6(in_reg_wire_3[190]),
    .out7(in_reg_wire_3[191])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_24
  (
    .sel(conf_out[1367:1344]),
    .in0(in_reg_wire_2[24]),
    .in1(in_reg_wire_2[56]),
    .in2(in_reg_wire_2[88]),
    .in3(in_reg_wire_2[120]),
    .in4(in_reg_wire_2[152]),
    .in5(in_reg_wire_2[184]),
    .in6(in_reg_wire_2[216]),
    .in7(in_reg_wire_2[248]),
    .out0(in_reg_wire_3[192]),
    .out1(in_reg_wire_3[193]),
    .out2(in_reg_wire_3[194]),
    .out3(in_reg_wire_3[195]),
    .out4(in_reg_wire_3[196]),
    .out5(in_reg_wire_3[197]),
    .out6(in_reg_wire_3[198]),
    .out7(in_reg_wire_3[199])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_25
  (
    .sel(conf_out[1391:1368]),
    .in0(in_reg_wire_2[25]),
    .in1(in_reg_wire_2[57]),
    .in2(in_reg_wire_2[89]),
    .in3(in_reg_wire_2[121]),
    .in4(in_reg_wire_2[153]),
    .in5(in_reg_wire_2[185]),
    .in6(in_reg_wire_2[217]),
    .in7(in_reg_wire_2[249]),
    .out0(in_reg_wire_3[200]),
    .out1(in_reg_wire_3[201]),
    .out2(in_reg_wire_3[202]),
    .out3(in_reg_wire_3[203]),
    .out4(in_reg_wire_3[204]),
    .out5(in_reg_wire_3[205]),
    .out6(in_reg_wire_3[206]),
    .out7(in_reg_wire_3[207])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_26
  (
    .sel(conf_out[1415:1392]),
    .in0(in_reg_wire_2[26]),
    .in1(in_reg_wire_2[58]),
    .in2(in_reg_wire_2[90]),
    .in3(in_reg_wire_2[122]),
    .in4(in_reg_wire_2[154]),
    .in5(in_reg_wire_2[186]),
    .in6(in_reg_wire_2[218]),
    .in7(in_reg_wire_2[250]),
    .out0(in_reg_wire_3[208]),
    .out1(in_reg_wire_3[209]),
    .out2(in_reg_wire_3[210]),
    .out3(in_reg_wire_3[211]),
    .out4(in_reg_wire_3[212]),
    .out5(in_reg_wire_3[213]),
    .out6(in_reg_wire_3[214]),
    .out7(in_reg_wire_3[215])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_27
  (
    .sel(conf_out[1439:1416]),
    .in0(in_reg_wire_2[27]),
    .in1(in_reg_wire_2[59]),
    .in2(in_reg_wire_2[91]),
    .in3(in_reg_wire_2[123]),
    .in4(in_reg_wire_2[155]),
    .in5(in_reg_wire_2[187]),
    .in6(in_reg_wire_2[219]),
    .in7(in_reg_wire_2[251]),
    .out0(in_reg_wire_3[216]),
    .out1(in_reg_wire_3[217]),
    .out2(in_reg_wire_3[218]),
    .out3(in_reg_wire_3[219]),
    .out4(in_reg_wire_3[220]),
    .out5(in_reg_wire_3[221]),
    .out6(in_reg_wire_3[222]),
    .out7(in_reg_wire_3[223])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_28
  (
    .sel(conf_out[1463:1440]),
    .in0(in_reg_wire_2[28]),
    .in1(in_reg_wire_2[60]),
    .in2(in_reg_wire_2[92]),
    .in3(in_reg_wire_2[124]),
    .in4(in_reg_wire_2[156]),
    .in5(in_reg_wire_2[188]),
    .in6(in_reg_wire_2[220]),
    .in7(in_reg_wire_2[252]),
    .out0(in_reg_wire_3[224]),
    .out1(in_reg_wire_3[225]),
    .out2(in_reg_wire_3[226]),
    .out3(in_reg_wire_3[227]),
    .out4(in_reg_wire_3[228]),
    .out5(in_reg_wire_3[229]),
    .out6(in_reg_wire_3[230]),
    .out7(in_reg_wire_3[231])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_29
  (
    .sel(conf_out[1487:1464]),
    .in0(in_reg_wire_2[29]),
    .in1(in_reg_wire_2[61]),
    .in2(in_reg_wire_2[93]),
    .in3(in_reg_wire_2[125]),
    .in4(in_reg_wire_2[157]),
    .in5(in_reg_wire_2[189]),
    .in6(in_reg_wire_2[221]),
    .in7(in_reg_wire_2[253]),
    .out0(in_reg_wire_3[232]),
    .out1(in_reg_wire_3[233]),
    .out2(in_reg_wire_3[234]),
    .out3(in_reg_wire_3[235]),
    .out4(in_reg_wire_3[236]),
    .out5(in_reg_wire_3[237]),
    .out6(in_reg_wire_3[238]),
    .out7(in_reg_wire_3[239])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_30
  (
    .sel(conf_out[1511:1488]),
    .in0(in_reg_wire_2[30]),
    .in1(in_reg_wire_2[62]),
    .in2(in_reg_wire_2[94]),
    .in3(in_reg_wire_2[126]),
    .in4(in_reg_wire_2[158]),
    .in5(in_reg_wire_2[190]),
    .in6(in_reg_wire_2[222]),
    .in7(in_reg_wire_2[254]),
    .out0(in_reg_wire_3[240]),
    .out1(in_reg_wire_3[241]),
    .out2(in_reg_wire_3[242]),
    .out3(in_reg_wire_3[243]),
    .out4(in_reg_wire_3[244]),
    .out5(in_reg_wire_3[245]),
    .out6(in_reg_wire_3[246]),
    .out7(in_reg_wire_3[247])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_31
  (
    .sel(conf_out[1535:1512]),
    .in0(in_reg_wire_2[31]),
    .in1(in_reg_wire_2[63]),
    .in2(in_reg_wire_2[95]),
    .in3(in_reg_wire_2[127]),
    .in4(in_reg_wire_2[159]),
    .in5(in_reg_wire_2[191]),
    .in6(in_reg_wire_2[223]),
    .in7(in_reg_wire_2[255]),
    .out0(in_reg_wire_3[248]),
    .out1(in_reg_wire_3[249]),
    .out2(in_reg_wire_3[250]),
    .out3(in_reg_wire_3[251]),
    .out4(in_reg_wire_3[252]),
    .out5(in_reg_wire_3[253]),
    .out6(in_reg_wire_3[254]),
    .out7(in_reg_wire_3[255])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_0
  (
    .sel(conf_out[1559:1536]),
    .in0(in_reg_wire_4[0]),
    .in1(in_reg_wire_4[32]),
    .in2(in_reg_wire_4[64]),
    .in3(in_reg_wire_4[96]),
    .in4(in_reg_wire_4[128]),
    .in5(in_reg_wire_4[160]),
    .in6(in_reg_wire_4[192]),
    .in7(in_reg_wire_4[224]),
    .out0(in_reg_wire_5[0]),
    .out1(in_reg_wire_5[1]),
    .out2(in_reg_wire_5[2]),
    .out3(in_reg_wire_5[3]),
    .out4(in_reg_wire_5[4]),
    .out5(in_reg_wire_5[5]),
    .out6(in_reg_wire_5[6]),
    .out7(in_reg_wire_5[7])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_1
  (
    .sel(conf_out[1583:1560]),
    .in0(in_reg_wire_4[1]),
    .in1(in_reg_wire_4[33]),
    .in2(in_reg_wire_4[65]),
    .in3(in_reg_wire_4[97]),
    .in4(in_reg_wire_4[129]),
    .in5(in_reg_wire_4[161]),
    .in6(in_reg_wire_4[193]),
    .in7(in_reg_wire_4[225]),
    .out0(in_reg_wire_5[8]),
    .out1(in_reg_wire_5[9]),
    .out2(in_reg_wire_5[10]),
    .out3(in_reg_wire_5[11]),
    .out4(in_reg_wire_5[12]),
    .out5(in_reg_wire_5[13]),
    .out6(in_reg_wire_5[14]),
    .out7(in_reg_wire_5[15])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_2
  (
    .sel(conf_out[1607:1584]),
    .in0(in_reg_wire_4[2]),
    .in1(in_reg_wire_4[34]),
    .in2(in_reg_wire_4[66]),
    .in3(in_reg_wire_4[98]),
    .in4(in_reg_wire_4[130]),
    .in5(in_reg_wire_4[162]),
    .in6(in_reg_wire_4[194]),
    .in7(in_reg_wire_4[226]),
    .out0(in_reg_wire_5[16]),
    .out1(in_reg_wire_5[17]),
    .out2(in_reg_wire_5[18]),
    .out3(in_reg_wire_5[19]),
    .out4(in_reg_wire_5[20]),
    .out5(in_reg_wire_5[21]),
    .out6(in_reg_wire_5[22]),
    .out7(in_reg_wire_5[23])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_3
  (
    .sel(conf_out[1631:1608]),
    .in0(in_reg_wire_4[3]),
    .in1(in_reg_wire_4[35]),
    .in2(in_reg_wire_4[67]),
    .in3(in_reg_wire_4[99]),
    .in4(in_reg_wire_4[131]),
    .in5(in_reg_wire_4[163]),
    .in6(in_reg_wire_4[195]),
    .in7(in_reg_wire_4[227]),
    .out0(in_reg_wire_5[24]),
    .out1(in_reg_wire_5[25]),
    .out2(in_reg_wire_5[26]),
    .out3(in_reg_wire_5[27]),
    .out4(in_reg_wire_5[28]),
    .out5(in_reg_wire_5[29]),
    .out6(in_reg_wire_5[30]),
    .out7(in_reg_wire_5[31])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_4
  (
    .sel(conf_out[1655:1632]),
    .in0(in_reg_wire_4[4]),
    .in1(in_reg_wire_4[36]),
    .in2(in_reg_wire_4[68]),
    .in3(in_reg_wire_4[100]),
    .in4(in_reg_wire_4[132]),
    .in5(in_reg_wire_4[164]),
    .in6(in_reg_wire_4[196]),
    .in7(in_reg_wire_4[228]),
    .out0(in_reg_wire_5[32]),
    .out1(in_reg_wire_5[33]),
    .out2(in_reg_wire_5[34]),
    .out3(in_reg_wire_5[35]),
    .out4(in_reg_wire_5[36]),
    .out5(in_reg_wire_5[37]),
    .out6(in_reg_wire_5[38]),
    .out7(in_reg_wire_5[39])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_5
  (
    .sel(conf_out[1679:1656]),
    .in0(in_reg_wire_4[5]),
    .in1(in_reg_wire_4[37]),
    .in2(in_reg_wire_4[69]),
    .in3(in_reg_wire_4[101]),
    .in4(in_reg_wire_4[133]),
    .in5(in_reg_wire_4[165]),
    .in6(in_reg_wire_4[197]),
    .in7(in_reg_wire_4[229]),
    .out0(in_reg_wire_5[40]),
    .out1(in_reg_wire_5[41]),
    .out2(in_reg_wire_5[42]),
    .out3(in_reg_wire_5[43]),
    .out4(in_reg_wire_5[44]),
    .out5(in_reg_wire_5[45]),
    .out6(in_reg_wire_5[46]),
    .out7(in_reg_wire_5[47])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_6
  (
    .sel(conf_out[1703:1680]),
    .in0(in_reg_wire_4[6]),
    .in1(in_reg_wire_4[38]),
    .in2(in_reg_wire_4[70]),
    .in3(in_reg_wire_4[102]),
    .in4(in_reg_wire_4[134]),
    .in5(in_reg_wire_4[166]),
    .in6(in_reg_wire_4[198]),
    .in7(in_reg_wire_4[230]),
    .out0(in_reg_wire_5[48]),
    .out1(in_reg_wire_5[49]),
    .out2(in_reg_wire_5[50]),
    .out3(in_reg_wire_5[51]),
    .out4(in_reg_wire_5[52]),
    .out5(in_reg_wire_5[53]),
    .out6(in_reg_wire_5[54]),
    .out7(in_reg_wire_5[55])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_7
  (
    .sel(conf_out[1727:1704]),
    .in0(in_reg_wire_4[7]),
    .in1(in_reg_wire_4[39]),
    .in2(in_reg_wire_4[71]),
    .in3(in_reg_wire_4[103]),
    .in4(in_reg_wire_4[135]),
    .in5(in_reg_wire_4[167]),
    .in6(in_reg_wire_4[199]),
    .in7(in_reg_wire_4[231]),
    .out0(in_reg_wire_5[56]),
    .out1(in_reg_wire_5[57]),
    .out2(in_reg_wire_5[58]),
    .out3(in_reg_wire_5[59]),
    .out4(in_reg_wire_5[60]),
    .out5(in_reg_wire_5[61]),
    .out6(in_reg_wire_5[62]),
    .out7(in_reg_wire_5[63])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_8
  (
    .sel(conf_out[1751:1728]),
    .in0(in_reg_wire_4[8]),
    .in1(in_reg_wire_4[40]),
    .in2(in_reg_wire_4[72]),
    .in3(in_reg_wire_4[104]),
    .in4(in_reg_wire_4[136]),
    .in5(in_reg_wire_4[168]),
    .in6(in_reg_wire_4[200]),
    .in7(in_reg_wire_4[232]),
    .out0(in_reg_wire_5[64]),
    .out1(in_reg_wire_5[65]),
    .out2(in_reg_wire_5[66]),
    .out3(in_reg_wire_5[67]),
    .out4(in_reg_wire_5[68]),
    .out5(in_reg_wire_5[69]),
    .out6(in_reg_wire_5[70]),
    .out7(in_reg_wire_5[71])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_9
  (
    .sel(conf_out[1775:1752]),
    .in0(in_reg_wire_4[9]),
    .in1(in_reg_wire_4[41]),
    .in2(in_reg_wire_4[73]),
    .in3(in_reg_wire_4[105]),
    .in4(in_reg_wire_4[137]),
    .in5(in_reg_wire_4[169]),
    .in6(in_reg_wire_4[201]),
    .in7(in_reg_wire_4[233]),
    .out0(in_reg_wire_5[72]),
    .out1(in_reg_wire_5[73]),
    .out2(in_reg_wire_5[74]),
    .out3(in_reg_wire_5[75]),
    .out4(in_reg_wire_5[76]),
    .out5(in_reg_wire_5[77]),
    .out6(in_reg_wire_5[78]),
    .out7(in_reg_wire_5[79])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_10
  (
    .sel(conf_out[1799:1776]),
    .in0(in_reg_wire_4[10]),
    .in1(in_reg_wire_4[42]),
    .in2(in_reg_wire_4[74]),
    .in3(in_reg_wire_4[106]),
    .in4(in_reg_wire_4[138]),
    .in5(in_reg_wire_4[170]),
    .in6(in_reg_wire_4[202]),
    .in7(in_reg_wire_4[234]),
    .out0(in_reg_wire_5[80]),
    .out1(in_reg_wire_5[81]),
    .out2(in_reg_wire_5[82]),
    .out3(in_reg_wire_5[83]),
    .out4(in_reg_wire_5[84]),
    .out5(in_reg_wire_5[85]),
    .out6(in_reg_wire_5[86]),
    .out7(in_reg_wire_5[87])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_11
  (
    .sel(conf_out[1823:1800]),
    .in0(in_reg_wire_4[11]),
    .in1(in_reg_wire_4[43]),
    .in2(in_reg_wire_4[75]),
    .in3(in_reg_wire_4[107]),
    .in4(in_reg_wire_4[139]),
    .in5(in_reg_wire_4[171]),
    .in6(in_reg_wire_4[203]),
    .in7(in_reg_wire_4[235]),
    .out0(in_reg_wire_5[88]),
    .out1(in_reg_wire_5[89]),
    .out2(in_reg_wire_5[90]),
    .out3(in_reg_wire_5[91]),
    .out4(in_reg_wire_5[92]),
    .out5(in_reg_wire_5[93]),
    .out6(in_reg_wire_5[94]),
    .out7(in_reg_wire_5[95])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_12
  (
    .sel(conf_out[1847:1824]),
    .in0(in_reg_wire_4[12]),
    .in1(in_reg_wire_4[44]),
    .in2(in_reg_wire_4[76]),
    .in3(in_reg_wire_4[108]),
    .in4(in_reg_wire_4[140]),
    .in5(in_reg_wire_4[172]),
    .in6(in_reg_wire_4[204]),
    .in7(in_reg_wire_4[236]),
    .out0(in_reg_wire_5[96]),
    .out1(in_reg_wire_5[97]),
    .out2(in_reg_wire_5[98]),
    .out3(in_reg_wire_5[99]),
    .out4(in_reg_wire_5[100]),
    .out5(in_reg_wire_5[101]),
    .out6(in_reg_wire_5[102]),
    .out7(in_reg_wire_5[103])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_13
  (
    .sel(conf_out[1871:1848]),
    .in0(in_reg_wire_4[13]),
    .in1(in_reg_wire_4[45]),
    .in2(in_reg_wire_4[77]),
    .in3(in_reg_wire_4[109]),
    .in4(in_reg_wire_4[141]),
    .in5(in_reg_wire_4[173]),
    .in6(in_reg_wire_4[205]),
    .in7(in_reg_wire_4[237]),
    .out0(in_reg_wire_5[104]),
    .out1(in_reg_wire_5[105]),
    .out2(in_reg_wire_5[106]),
    .out3(in_reg_wire_5[107]),
    .out4(in_reg_wire_5[108]),
    .out5(in_reg_wire_5[109]),
    .out6(in_reg_wire_5[110]),
    .out7(in_reg_wire_5[111])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_14
  (
    .sel(conf_out[1895:1872]),
    .in0(in_reg_wire_4[14]),
    .in1(in_reg_wire_4[46]),
    .in2(in_reg_wire_4[78]),
    .in3(in_reg_wire_4[110]),
    .in4(in_reg_wire_4[142]),
    .in5(in_reg_wire_4[174]),
    .in6(in_reg_wire_4[206]),
    .in7(in_reg_wire_4[238]),
    .out0(in_reg_wire_5[112]),
    .out1(in_reg_wire_5[113]),
    .out2(in_reg_wire_5[114]),
    .out3(in_reg_wire_5[115]),
    .out4(in_reg_wire_5[116]),
    .out5(in_reg_wire_5[117]),
    .out6(in_reg_wire_5[118]),
    .out7(in_reg_wire_5[119])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_15
  (
    .sel(conf_out[1919:1896]),
    .in0(in_reg_wire_4[15]),
    .in1(in_reg_wire_4[47]),
    .in2(in_reg_wire_4[79]),
    .in3(in_reg_wire_4[111]),
    .in4(in_reg_wire_4[143]),
    .in5(in_reg_wire_4[175]),
    .in6(in_reg_wire_4[207]),
    .in7(in_reg_wire_4[239]),
    .out0(in_reg_wire_5[120]),
    .out1(in_reg_wire_5[121]),
    .out2(in_reg_wire_5[122]),
    .out3(in_reg_wire_5[123]),
    .out4(in_reg_wire_5[124]),
    .out5(in_reg_wire_5[125]),
    .out6(in_reg_wire_5[126]),
    .out7(in_reg_wire_5[127])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_16
  (
    .sel(conf_out[1943:1920]),
    .in0(in_reg_wire_4[16]),
    .in1(in_reg_wire_4[48]),
    .in2(in_reg_wire_4[80]),
    .in3(in_reg_wire_4[112]),
    .in4(in_reg_wire_4[144]),
    .in5(in_reg_wire_4[176]),
    .in6(in_reg_wire_4[208]),
    .in7(in_reg_wire_4[240]),
    .out0(in_reg_wire_5[128]),
    .out1(in_reg_wire_5[129]),
    .out2(in_reg_wire_5[130]),
    .out3(in_reg_wire_5[131]),
    .out4(in_reg_wire_5[132]),
    .out5(in_reg_wire_5[133]),
    .out6(in_reg_wire_5[134]),
    .out7(in_reg_wire_5[135])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_17
  (
    .sel(conf_out[1967:1944]),
    .in0(in_reg_wire_4[17]),
    .in1(in_reg_wire_4[49]),
    .in2(in_reg_wire_4[81]),
    .in3(in_reg_wire_4[113]),
    .in4(in_reg_wire_4[145]),
    .in5(in_reg_wire_4[177]),
    .in6(in_reg_wire_4[209]),
    .in7(in_reg_wire_4[241]),
    .out0(in_reg_wire_5[136]),
    .out1(in_reg_wire_5[137]),
    .out2(in_reg_wire_5[138]),
    .out3(in_reg_wire_5[139]),
    .out4(in_reg_wire_5[140]),
    .out5(in_reg_wire_5[141]),
    .out6(in_reg_wire_5[142]),
    .out7(in_reg_wire_5[143])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_18
  (
    .sel(conf_out[1991:1968]),
    .in0(in_reg_wire_4[18]),
    .in1(in_reg_wire_4[50]),
    .in2(in_reg_wire_4[82]),
    .in3(in_reg_wire_4[114]),
    .in4(in_reg_wire_4[146]),
    .in5(in_reg_wire_4[178]),
    .in6(in_reg_wire_4[210]),
    .in7(in_reg_wire_4[242]),
    .out0(in_reg_wire_5[144]),
    .out1(in_reg_wire_5[145]),
    .out2(in_reg_wire_5[146]),
    .out3(in_reg_wire_5[147]),
    .out4(in_reg_wire_5[148]),
    .out5(in_reg_wire_5[149]),
    .out6(in_reg_wire_5[150]),
    .out7(in_reg_wire_5[151])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_19
  (
    .sel(conf_out[2015:1992]),
    .in0(in_reg_wire_4[19]),
    .in1(in_reg_wire_4[51]),
    .in2(in_reg_wire_4[83]),
    .in3(in_reg_wire_4[115]),
    .in4(in_reg_wire_4[147]),
    .in5(in_reg_wire_4[179]),
    .in6(in_reg_wire_4[211]),
    .in7(in_reg_wire_4[243]),
    .out0(in_reg_wire_5[152]),
    .out1(in_reg_wire_5[153]),
    .out2(in_reg_wire_5[154]),
    .out3(in_reg_wire_5[155]),
    .out4(in_reg_wire_5[156]),
    .out5(in_reg_wire_5[157]),
    .out6(in_reg_wire_5[158]),
    .out7(in_reg_wire_5[159])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_20
  (
    .sel(conf_out[2039:2016]),
    .in0(in_reg_wire_4[20]),
    .in1(in_reg_wire_4[52]),
    .in2(in_reg_wire_4[84]),
    .in3(in_reg_wire_4[116]),
    .in4(in_reg_wire_4[148]),
    .in5(in_reg_wire_4[180]),
    .in6(in_reg_wire_4[212]),
    .in7(in_reg_wire_4[244]),
    .out0(in_reg_wire_5[160]),
    .out1(in_reg_wire_5[161]),
    .out2(in_reg_wire_5[162]),
    .out3(in_reg_wire_5[163]),
    .out4(in_reg_wire_5[164]),
    .out5(in_reg_wire_5[165]),
    .out6(in_reg_wire_5[166]),
    .out7(in_reg_wire_5[167])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_21
  (
    .sel(conf_out[2063:2040]),
    .in0(in_reg_wire_4[21]),
    .in1(in_reg_wire_4[53]),
    .in2(in_reg_wire_4[85]),
    .in3(in_reg_wire_4[117]),
    .in4(in_reg_wire_4[149]),
    .in5(in_reg_wire_4[181]),
    .in6(in_reg_wire_4[213]),
    .in7(in_reg_wire_4[245]),
    .out0(in_reg_wire_5[168]),
    .out1(in_reg_wire_5[169]),
    .out2(in_reg_wire_5[170]),
    .out3(in_reg_wire_5[171]),
    .out4(in_reg_wire_5[172]),
    .out5(in_reg_wire_5[173]),
    .out6(in_reg_wire_5[174]),
    .out7(in_reg_wire_5[175])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_22
  (
    .sel(conf_out[2087:2064]),
    .in0(in_reg_wire_4[22]),
    .in1(in_reg_wire_4[54]),
    .in2(in_reg_wire_4[86]),
    .in3(in_reg_wire_4[118]),
    .in4(in_reg_wire_4[150]),
    .in5(in_reg_wire_4[182]),
    .in6(in_reg_wire_4[214]),
    .in7(in_reg_wire_4[246]),
    .out0(in_reg_wire_5[176]),
    .out1(in_reg_wire_5[177]),
    .out2(in_reg_wire_5[178]),
    .out3(in_reg_wire_5[179]),
    .out4(in_reg_wire_5[180]),
    .out5(in_reg_wire_5[181]),
    .out6(in_reg_wire_5[182]),
    .out7(in_reg_wire_5[183])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_23
  (
    .sel(conf_out[2111:2088]),
    .in0(in_reg_wire_4[23]),
    .in1(in_reg_wire_4[55]),
    .in2(in_reg_wire_4[87]),
    .in3(in_reg_wire_4[119]),
    .in4(in_reg_wire_4[151]),
    .in5(in_reg_wire_4[183]),
    .in6(in_reg_wire_4[215]),
    .in7(in_reg_wire_4[247]),
    .out0(in_reg_wire_5[184]),
    .out1(in_reg_wire_5[185]),
    .out2(in_reg_wire_5[186]),
    .out3(in_reg_wire_5[187]),
    .out4(in_reg_wire_5[188]),
    .out5(in_reg_wire_5[189]),
    .out6(in_reg_wire_5[190]),
    .out7(in_reg_wire_5[191])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_24
  (
    .sel(conf_out[2135:2112]),
    .in0(in_reg_wire_4[24]),
    .in1(in_reg_wire_4[56]),
    .in2(in_reg_wire_4[88]),
    .in3(in_reg_wire_4[120]),
    .in4(in_reg_wire_4[152]),
    .in5(in_reg_wire_4[184]),
    .in6(in_reg_wire_4[216]),
    .in7(in_reg_wire_4[248]),
    .out0(in_reg_wire_5[192]),
    .out1(in_reg_wire_5[193]),
    .out2(in_reg_wire_5[194]),
    .out3(in_reg_wire_5[195]),
    .out4(in_reg_wire_5[196]),
    .out5(in_reg_wire_5[197]),
    .out6(in_reg_wire_5[198]),
    .out7(in_reg_wire_5[199])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_25
  (
    .sel(conf_out[2159:2136]),
    .in0(in_reg_wire_4[25]),
    .in1(in_reg_wire_4[57]),
    .in2(in_reg_wire_4[89]),
    .in3(in_reg_wire_4[121]),
    .in4(in_reg_wire_4[153]),
    .in5(in_reg_wire_4[185]),
    .in6(in_reg_wire_4[217]),
    .in7(in_reg_wire_4[249]),
    .out0(in_reg_wire_5[200]),
    .out1(in_reg_wire_5[201]),
    .out2(in_reg_wire_5[202]),
    .out3(in_reg_wire_5[203]),
    .out4(in_reg_wire_5[204]),
    .out5(in_reg_wire_5[205]),
    .out6(in_reg_wire_5[206]),
    .out7(in_reg_wire_5[207])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_26
  (
    .sel(conf_out[2183:2160]),
    .in0(in_reg_wire_4[26]),
    .in1(in_reg_wire_4[58]),
    .in2(in_reg_wire_4[90]),
    .in3(in_reg_wire_4[122]),
    .in4(in_reg_wire_4[154]),
    .in5(in_reg_wire_4[186]),
    .in6(in_reg_wire_4[218]),
    .in7(in_reg_wire_4[250]),
    .out0(in_reg_wire_5[208]),
    .out1(in_reg_wire_5[209]),
    .out2(in_reg_wire_5[210]),
    .out3(in_reg_wire_5[211]),
    .out4(in_reg_wire_5[212]),
    .out5(in_reg_wire_5[213]),
    .out6(in_reg_wire_5[214]),
    .out7(in_reg_wire_5[215])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_27
  (
    .sel(conf_out[2207:2184]),
    .in0(in_reg_wire_4[27]),
    .in1(in_reg_wire_4[59]),
    .in2(in_reg_wire_4[91]),
    .in3(in_reg_wire_4[123]),
    .in4(in_reg_wire_4[155]),
    .in5(in_reg_wire_4[187]),
    .in6(in_reg_wire_4[219]),
    .in7(in_reg_wire_4[251]),
    .out0(in_reg_wire_5[216]),
    .out1(in_reg_wire_5[217]),
    .out2(in_reg_wire_5[218]),
    .out3(in_reg_wire_5[219]),
    .out4(in_reg_wire_5[220]),
    .out5(in_reg_wire_5[221]),
    .out6(in_reg_wire_5[222]),
    .out7(in_reg_wire_5[223])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_28
  (
    .sel(conf_out[2231:2208]),
    .in0(in_reg_wire_4[28]),
    .in1(in_reg_wire_4[60]),
    .in2(in_reg_wire_4[92]),
    .in3(in_reg_wire_4[124]),
    .in4(in_reg_wire_4[156]),
    .in5(in_reg_wire_4[188]),
    .in6(in_reg_wire_4[220]),
    .in7(in_reg_wire_4[252]),
    .out0(in_reg_wire_5[224]),
    .out1(in_reg_wire_5[225]),
    .out2(in_reg_wire_5[226]),
    .out3(in_reg_wire_5[227]),
    .out4(in_reg_wire_5[228]),
    .out5(in_reg_wire_5[229]),
    .out6(in_reg_wire_5[230]),
    .out7(in_reg_wire_5[231])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_29
  (
    .sel(conf_out[2255:2232]),
    .in0(in_reg_wire_4[29]),
    .in1(in_reg_wire_4[61]),
    .in2(in_reg_wire_4[93]),
    .in3(in_reg_wire_4[125]),
    .in4(in_reg_wire_4[157]),
    .in5(in_reg_wire_4[189]),
    .in6(in_reg_wire_4[221]),
    .in7(in_reg_wire_4[253]),
    .out0(in_reg_wire_5[232]),
    .out1(in_reg_wire_5[233]),
    .out2(in_reg_wire_5[234]),
    .out3(in_reg_wire_5[235]),
    .out4(in_reg_wire_5[236]),
    .out5(in_reg_wire_5[237]),
    .out6(in_reg_wire_5[238]),
    .out7(in_reg_wire_5[239])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_30
  (
    .sel(conf_out[2279:2256]),
    .in0(in_reg_wire_4[30]),
    .in1(in_reg_wire_4[62]),
    .in2(in_reg_wire_4[94]),
    .in3(in_reg_wire_4[126]),
    .in4(in_reg_wire_4[158]),
    .in5(in_reg_wire_4[190]),
    .in6(in_reg_wire_4[222]),
    .in7(in_reg_wire_4[254]),
    .out0(in_reg_wire_5[240]),
    .out1(in_reg_wire_5[241]),
    .out2(in_reg_wire_5[242]),
    .out3(in_reg_wire_5[243]),
    .out4(in_reg_wire_5[244]),
    .out5(in_reg_wire_5[245]),
    .out6(in_reg_wire_5[246]),
    .out7(in_reg_wire_5[247])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_31
  (
    .sel(conf_out[2303:2280]),
    .in0(in_reg_wire_4[31]),
    .in1(in_reg_wire_4[63]),
    .in2(in_reg_wire_4[95]),
    .in3(in_reg_wire_4[127]),
    .in4(in_reg_wire_4[159]),
    .in5(in_reg_wire_4[191]),
    .in6(in_reg_wire_4[223]),
    .in7(in_reg_wire_4[255]),
    .out0(in_reg_wire_5[248]),
    .out1(in_reg_wire_5[249]),
    .out2(in_reg_wire_5[250]),
    .out3(in_reg_wire_5[251]),
    .out4(in_reg_wire_5[252]),
    .out5(in_reg_wire_5[253]),
    .out6(in_reg_wire_5[254]),
    .out7(in_reg_wire_5[255])
  );

endmodule