module cgra0_top
(
  input clk,
  input rst,
  input en,
  input [64-1:0] conf_bus_in,
  output [8-1:0] fifo_in_re,
  input [128-1:0] fifo_in_data,
  output [8-1:0] fifo_out_we,
  output [128-1:0] fifo_out_data
);


  wire [64-1:0] conf_bus [0:130-1];
  wire [16-1:0] pe2neta [0:128-1];
  wire [16-1:0] pe2netb [0:128-1];
  wire [16-1:0] net2pea [0:128-1];
  wire [16-1:0] net2peb [0:128-1];
  wire [128-1:0] pe2net_branch;
  wire [128-1:0] net_branch2peb;


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  reg_conf_bus_in2
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus_in),
    .out(conf_bus[0])
  );


  cgra0_pe_in
  #(
    .PE_ID(1)
  )
  pe_io_in_1
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[0]),
    .branch_in(net_branch2peb[0]),
    .branch_out(pe2net_branch[0]),
    .fifo_re(fifo_in_re[0]),
    .fifo_data(fifo_in_data[15:0]),
    .ina(net2pea[0]),
    .inb(net2peb[0]),
    .outa(pe2neta[0]),
    .outb(pe2netb[0])
  );


  cgra0_pe_in
  #(
    .PE_ID(2)
  )
  pe_io_in_2
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[1]),
    .branch_in(net_branch2peb[1]),
    .branch_out(pe2net_branch[1]),
    .fifo_re(fifo_in_re[1]),
    .fifo_data(fifo_in_data[31:16]),
    .ina(net2pea[1]),
    .inb(net2peb[1]),
    .outa(pe2neta[1]),
    .outb(pe2netb[1])
  );


  cgra0_pe_in
  #(
    .PE_ID(3)
  )
  pe_io_in_3
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[2]),
    .branch_in(net_branch2peb[2]),
    .branch_out(pe2net_branch[2]),
    .fifo_re(fifo_in_re[2]),
    .fifo_data(fifo_in_data[47:32]),
    .ina(net2pea[2]),
    .inb(net2peb[2]),
    .outa(pe2neta[2]),
    .outb(pe2netb[2])
  );


  cgra0_pe_in
  #(
    .PE_ID(4)
  )
  pe_io_in_4
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[3]),
    .branch_in(net_branch2peb[3]),
    .branch_out(pe2net_branch[3]),
    .fifo_re(fifo_in_re[3]),
    .fifo_data(fifo_in_data[63:48]),
    .ina(net2pea[3]),
    .inb(net2peb[3]),
    .outa(pe2neta[3]),
    .outb(pe2netb[3])
  );


  cgra0_pe_in
  #(
    .PE_ID(5)
  )
  pe_io_in_5
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[4]),
    .branch_in(net_branch2peb[4]),
    .branch_out(pe2net_branch[4]),
    .fifo_re(fifo_in_re[4]),
    .fifo_data(fifo_in_data[79:64]),
    .ina(net2pea[4]),
    .inb(net2peb[4]),
    .outa(pe2neta[4]),
    .outb(pe2netb[4])
  );


  cgra0_pe_in
  #(
    .PE_ID(6)
  )
  pe_io_in_6
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[5]),
    .branch_in(net_branch2peb[5]),
    .branch_out(pe2net_branch[5]),
    .fifo_re(fifo_in_re[5]),
    .fifo_data(fifo_in_data[95:80]),
    .ina(net2pea[5]),
    .inb(net2peb[5]),
    .outa(pe2neta[5]),
    .outb(pe2netb[5])
  );


  cgra0_pe_in
  #(
    .PE_ID(7)
  )
  pe_io_in_7
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[6]),
    .branch_in(net_branch2peb[6]),
    .branch_out(pe2net_branch[6]),
    .fifo_re(fifo_in_re[6]),
    .fifo_data(fifo_in_data[111:96]),
    .ina(net2pea[6]),
    .inb(net2peb[6]),
    .outa(pe2neta[6]),
    .outb(pe2netb[6])
  );


  cgra0_pe_in
  #(
    .PE_ID(8)
  )
  pe_io_in_8
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[7]),
    .branch_in(net_branch2peb[7]),
    .branch_out(pe2net_branch[7]),
    .fifo_re(fifo_in_re[7]),
    .fifo_data(fifo_in_data[127:112]),
    .ina(net2pea[7]),
    .inb(net2peb[7]),
    .outa(pe2neta[7]),
    .outb(pe2netb[7])
  );


  cgra0_pe
  #(
    .PE_ID(9)
  )
  pe_9
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[8]),
    .branch_in(net_branch2peb[8]),
    .branch_out(pe2net_branch[8]),
    .ina(net2pea[8]),
    .inb(net2peb[8]),
    .outa(pe2neta[8]),
    .outb(pe2netb[8])
  );


  cgra0_pe
  #(
    .PE_ID(10)
  )
  pe_10
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[9]),
    .branch_in(net_branch2peb[9]),
    .branch_out(pe2net_branch[9]),
    .ina(net2pea[9]),
    .inb(net2peb[9]),
    .outa(pe2neta[9]),
    .outb(pe2netb[9])
  );


  cgra0_pe
  #(
    .PE_ID(11)
  )
  pe_11
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[10]),
    .branch_in(net_branch2peb[10]),
    .branch_out(pe2net_branch[10]),
    .ina(net2pea[10]),
    .inb(net2peb[10]),
    .outa(pe2neta[10]),
    .outb(pe2netb[10])
  );


  cgra0_pe
  #(
    .PE_ID(12)
  )
  pe_12
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[11]),
    .branch_in(net_branch2peb[11]),
    .branch_out(pe2net_branch[11]),
    .ina(net2pea[11]),
    .inb(net2peb[11]),
    .outa(pe2neta[11]),
    .outb(pe2netb[11])
  );


  cgra0_pe
  #(
    .PE_ID(13)
  )
  pe_13
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[12]),
    .branch_in(net_branch2peb[12]),
    .branch_out(pe2net_branch[12]),
    .ina(net2pea[12]),
    .inb(net2peb[12]),
    .outa(pe2neta[12]),
    .outb(pe2netb[12])
  );


  cgra0_pe
  #(
    .PE_ID(14)
  )
  pe_14
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[13]),
    .branch_in(net_branch2peb[13]),
    .branch_out(pe2net_branch[13]),
    .ina(net2pea[13]),
    .inb(net2peb[13]),
    .outa(pe2neta[13]),
    .outb(pe2netb[13])
  );


  cgra0_pe
  #(
    .PE_ID(15)
  )
  pe_15
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[14]),
    .branch_in(net_branch2peb[14]),
    .branch_out(pe2net_branch[14]),
    .ina(net2pea[14]),
    .inb(net2peb[14]),
    .outa(pe2neta[14]),
    .outb(pe2netb[14])
  );


  cgra0_pe
  #(
    .PE_ID(16)
  )
  pe_16
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[15]),
    .branch_in(net_branch2peb[15]),
    .branch_out(pe2net_branch[15]),
    .ina(net2pea[15]),
    .inb(net2peb[15]),
    .outa(pe2neta[15]),
    .outb(pe2netb[15])
  );


  cgra0_pe
  #(
    .PE_ID(17)
  )
  pe_17
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[16]),
    .branch_in(net_branch2peb[16]),
    .branch_out(pe2net_branch[16]),
    .ina(net2pea[16]),
    .inb(net2peb[16]),
    .outa(pe2neta[16]),
    .outb(pe2netb[16])
  );


  cgra0_pe
  #(
    .PE_ID(18)
  )
  pe_18
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[17]),
    .branch_in(net_branch2peb[17]),
    .branch_out(pe2net_branch[17]),
    .ina(net2pea[17]),
    .inb(net2peb[17]),
    .outa(pe2neta[17]),
    .outb(pe2netb[17])
  );


  cgra0_pe
  #(
    .PE_ID(19)
  )
  pe_19
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[18]),
    .branch_in(net_branch2peb[18]),
    .branch_out(pe2net_branch[18]),
    .ina(net2pea[18]),
    .inb(net2peb[18]),
    .outa(pe2neta[18]),
    .outb(pe2netb[18])
  );


  cgra0_pe
  #(
    .PE_ID(20)
  )
  pe_20
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[19]),
    .branch_in(net_branch2peb[19]),
    .branch_out(pe2net_branch[19]),
    .ina(net2pea[19]),
    .inb(net2peb[19]),
    .outa(pe2neta[19]),
    .outb(pe2netb[19])
  );


  cgra0_pe
  #(
    .PE_ID(21)
  )
  pe_21
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[20]),
    .branch_in(net_branch2peb[20]),
    .branch_out(pe2net_branch[20]),
    .ina(net2pea[20]),
    .inb(net2peb[20]),
    .outa(pe2neta[20]),
    .outb(pe2netb[20])
  );


  cgra0_pe
  #(
    .PE_ID(22)
  )
  pe_22
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[21]),
    .branch_in(net_branch2peb[21]),
    .branch_out(pe2net_branch[21]),
    .ina(net2pea[21]),
    .inb(net2peb[21]),
    .outa(pe2neta[21]),
    .outb(pe2netb[21])
  );


  cgra0_pe
  #(
    .PE_ID(23)
  )
  pe_23
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[22]),
    .branch_in(net_branch2peb[22]),
    .branch_out(pe2net_branch[22]),
    .ina(net2pea[22]),
    .inb(net2peb[22]),
    .outa(pe2neta[22]),
    .outb(pe2netb[22])
  );


  cgra0_pe
  #(
    .PE_ID(24)
  )
  pe_24
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[23]),
    .branch_in(net_branch2peb[23]),
    .branch_out(pe2net_branch[23]),
    .ina(net2pea[23]),
    .inb(net2peb[23]),
    .outa(pe2neta[23]),
    .outb(pe2netb[23])
  );


  cgra0_pe
  #(
    .PE_ID(25)
  )
  pe_25
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[24]),
    .branch_in(net_branch2peb[24]),
    .branch_out(pe2net_branch[24]),
    .ina(net2pea[24]),
    .inb(net2peb[24]),
    .outa(pe2neta[24]),
    .outb(pe2netb[24])
  );


  cgra0_pe
  #(
    .PE_ID(26)
  )
  pe_26
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[25]),
    .branch_in(net_branch2peb[25]),
    .branch_out(pe2net_branch[25]),
    .ina(net2pea[25]),
    .inb(net2peb[25]),
    .outa(pe2neta[25]),
    .outb(pe2netb[25])
  );


  cgra0_pe
  #(
    .PE_ID(27)
  )
  pe_27
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[26]),
    .branch_in(net_branch2peb[26]),
    .branch_out(pe2net_branch[26]),
    .ina(net2pea[26]),
    .inb(net2peb[26]),
    .outa(pe2neta[26]),
    .outb(pe2netb[26])
  );


  cgra0_pe
  #(
    .PE_ID(28)
  )
  pe_28
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[27]),
    .branch_in(net_branch2peb[27]),
    .branch_out(pe2net_branch[27]),
    .ina(net2pea[27]),
    .inb(net2peb[27]),
    .outa(pe2neta[27]),
    .outb(pe2netb[27])
  );


  cgra0_pe
  #(
    .PE_ID(29)
  )
  pe_29
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[28]),
    .branch_in(net_branch2peb[28]),
    .branch_out(pe2net_branch[28]),
    .ina(net2pea[28]),
    .inb(net2peb[28]),
    .outa(pe2neta[28]),
    .outb(pe2netb[28])
  );


  cgra0_pe
  #(
    .PE_ID(30)
  )
  pe_30
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[29]),
    .branch_in(net_branch2peb[29]),
    .branch_out(pe2net_branch[29]),
    .ina(net2pea[29]),
    .inb(net2peb[29]),
    .outa(pe2neta[29]),
    .outb(pe2netb[29])
  );


  cgra0_pe
  #(
    .PE_ID(31)
  )
  pe_31
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[30]),
    .branch_in(net_branch2peb[30]),
    .branch_out(pe2net_branch[30]),
    .ina(net2pea[30]),
    .inb(net2peb[30]),
    .outa(pe2neta[30]),
    .outb(pe2netb[30])
  );


  cgra0_pe
  #(
    .PE_ID(32)
  )
  pe_32
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[31]),
    .branch_in(net_branch2peb[31]),
    .branch_out(pe2net_branch[31]),
    .ina(net2pea[31]),
    .inb(net2peb[31]),
    .outa(pe2neta[31]),
    .outb(pe2netb[31])
  );


  cgra0_pe
  #(
    .PE_ID(33)
  )
  pe_33
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[32]),
    .branch_in(net_branch2peb[32]),
    .branch_out(pe2net_branch[32]),
    .ina(net2pea[32]),
    .inb(net2peb[32]),
    .outa(pe2neta[32]),
    .outb(pe2netb[32])
  );


  cgra0_pe
  #(
    .PE_ID(34)
  )
  pe_34
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[33]),
    .branch_in(net_branch2peb[33]),
    .branch_out(pe2net_branch[33]),
    .ina(net2pea[33]),
    .inb(net2peb[33]),
    .outa(pe2neta[33]),
    .outb(pe2netb[33])
  );


  cgra0_pe
  #(
    .PE_ID(35)
  )
  pe_35
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[34]),
    .branch_in(net_branch2peb[34]),
    .branch_out(pe2net_branch[34]),
    .ina(net2pea[34]),
    .inb(net2peb[34]),
    .outa(pe2neta[34]),
    .outb(pe2netb[34])
  );


  cgra0_pe
  #(
    .PE_ID(36)
  )
  pe_36
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[35]),
    .branch_in(net_branch2peb[35]),
    .branch_out(pe2net_branch[35]),
    .ina(net2pea[35]),
    .inb(net2peb[35]),
    .outa(pe2neta[35]),
    .outb(pe2netb[35])
  );


  cgra0_pe
  #(
    .PE_ID(37)
  )
  pe_37
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[36]),
    .branch_in(net_branch2peb[36]),
    .branch_out(pe2net_branch[36]),
    .ina(net2pea[36]),
    .inb(net2peb[36]),
    .outa(pe2neta[36]),
    .outb(pe2netb[36])
  );


  cgra0_pe
  #(
    .PE_ID(38)
  )
  pe_38
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[37]),
    .branch_in(net_branch2peb[37]),
    .branch_out(pe2net_branch[37]),
    .ina(net2pea[37]),
    .inb(net2peb[37]),
    .outa(pe2neta[37]),
    .outb(pe2netb[37])
  );


  cgra0_pe
  #(
    .PE_ID(39)
  )
  pe_39
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[38]),
    .branch_in(net_branch2peb[38]),
    .branch_out(pe2net_branch[38]),
    .ina(net2pea[38]),
    .inb(net2peb[38]),
    .outa(pe2neta[38]),
    .outb(pe2netb[38])
  );


  cgra0_pe
  #(
    .PE_ID(40)
  )
  pe_40
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[39]),
    .branch_in(net_branch2peb[39]),
    .branch_out(pe2net_branch[39]),
    .ina(net2pea[39]),
    .inb(net2peb[39]),
    .outa(pe2neta[39]),
    .outb(pe2netb[39])
  );


  cgra0_pe
  #(
    .PE_ID(41)
  )
  pe_41
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[40]),
    .branch_in(net_branch2peb[40]),
    .branch_out(pe2net_branch[40]),
    .ina(net2pea[40]),
    .inb(net2peb[40]),
    .outa(pe2neta[40]),
    .outb(pe2netb[40])
  );


  cgra0_pe
  #(
    .PE_ID(42)
  )
  pe_42
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[41]),
    .branch_in(net_branch2peb[41]),
    .branch_out(pe2net_branch[41]),
    .ina(net2pea[41]),
    .inb(net2peb[41]),
    .outa(pe2neta[41]),
    .outb(pe2netb[41])
  );


  cgra0_pe
  #(
    .PE_ID(43)
  )
  pe_43
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[42]),
    .branch_in(net_branch2peb[42]),
    .branch_out(pe2net_branch[42]),
    .ina(net2pea[42]),
    .inb(net2peb[42]),
    .outa(pe2neta[42]),
    .outb(pe2netb[42])
  );


  cgra0_pe
  #(
    .PE_ID(44)
  )
  pe_44
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[43]),
    .branch_in(net_branch2peb[43]),
    .branch_out(pe2net_branch[43]),
    .ina(net2pea[43]),
    .inb(net2peb[43]),
    .outa(pe2neta[43]),
    .outb(pe2netb[43])
  );


  cgra0_pe
  #(
    .PE_ID(45)
  )
  pe_45
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[44]),
    .branch_in(net_branch2peb[44]),
    .branch_out(pe2net_branch[44]),
    .ina(net2pea[44]),
    .inb(net2peb[44]),
    .outa(pe2neta[44]),
    .outb(pe2netb[44])
  );


  cgra0_pe
  #(
    .PE_ID(46)
  )
  pe_46
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[45]),
    .branch_in(net_branch2peb[45]),
    .branch_out(pe2net_branch[45]),
    .ina(net2pea[45]),
    .inb(net2peb[45]),
    .outa(pe2neta[45]),
    .outb(pe2netb[45])
  );


  cgra0_pe
  #(
    .PE_ID(47)
  )
  pe_47
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[46]),
    .branch_in(net_branch2peb[46]),
    .branch_out(pe2net_branch[46]),
    .ina(net2pea[46]),
    .inb(net2peb[46]),
    .outa(pe2neta[46]),
    .outb(pe2netb[46])
  );


  cgra0_pe
  #(
    .PE_ID(48)
  )
  pe_48
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[47]),
    .branch_in(net_branch2peb[47]),
    .branch_out(pe2net_branch[47]),
    .ina(net2pea[47]),
    .inb(net2peb[47]),
    .outa(pe2neta[47]),
    .outb(pe2netb[47])
  );


  cgra0_pe
  #(
    .PE_ID(49)
  )
  pe_49
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[48]),
    .branch_in(net_branch2peb[48]),
    .branch_out(pe2net_branch[48]),
    .ina(net2pea[48]),
    .inb(net2peb[48]),
    .outa(pe2neta[48]),
    .outb(pe2netb[48])
  );


  cgra0_pe
  #(
    .PE_ID(50)
  )
  pe_50
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[49]),
    .branch_in(net_branch2peb[49]),
    .branch_out(pe2net_branch[49]),
    .ina(net2pea[49]),
    .inb(net2peb[49]),
    .outa(pe2neta[49]),
    .outb(pe2netb[49])
  );


  cgra0_pe
  #(
    .PE_ID(51)
  )
  pe_51
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[50]),
    .branch_in(net_branch2peb[50]),
    .branch_out(pe2net_branch[50]),
    .ina(net2pea[50]),
    .inb(net2peb[50]),
    .outa(pe2neta[50]),
    .outb(pe2netb[50])
  );


  cgra0_pe
  #(
    .PE_ID(52)
  )
  pe_52
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[51]),
    .branch_in(net_branch2peb[51]),
    .branch_out(pe2net_branch[51]),
    .ina(net2pea[51]),
    .inb(net2peb[51]),
    .outa(pe2neta[51]),
    .outb(pe2netb[51])
  );


  cgra0_pe
  #(
    .PE_ID(53)
  )
  pe_53
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[52]),
    .branch_in(net_branch2peb[52]),
    .branch_out(pe2net_branch[52]),
    .ina(net2pea[52]),
    .inb(net2peb[52]),
    .outa(pe2neta[52]),
    .outb(pe2netb[52])
  );


  cgra0_pe
  #(
    .PE_ID(54)
  )
  pe_54
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[53]),
    .branch_in(net_branch2peb[53]),
    .branch_out(pe2net_branch[53]),
    .ina(net2pea[53]),
    .inb(net2peb[53]),
    .outa(pe2neta[53]),
    .outb(pe2netb[53])
  );


  cgra0_pe
  #(
    .PE_ID(55)
  )
  pe_55
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[54]),
    .branch_in(net_branch2peb[54]),
    .branch_out(pe2net_branch[54]),
    .ina(net2pea[54]),
    .inb(net2peb[54]),
    .outa(pe2neta[54]),
    .outb(pe2netb[54])
  );


  cgra0_pe
  #(
    .PE_ID(56)
  )
  pe_56
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[55]),
    .branch_in(net_branch2peb[55]),
    .branch_out(pe2net_branch[55]),
    .ina(net2pea[55]),
    .inb(net2peb[55]),
    .outa(pe2neta[55]),
    .outb(pe2netb[55])
  );


  cgra0_pe
  #(
    .PE_ID(57)
  )
  pe_57
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[56]),
    .branch_in(net_branch2peb[56]),
    .branch_out(pe2net_branch[56]),
    .ina(net2pea[56]),
    .inb(net2peb[56]),
    .outa(pe2neta[56]),
    .outb(pe2netb[56])
  );


  cgra0_pe
  #(
    .PE_ID(58)
  )
  pe_58
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[57]),
    .branch_in(net_branch2peb[57]),
    .branch_out(pe2net_branch[57]),
    .ina(net2pea[57]),
    .inb(net2peb[57]),
    .outa(pe2neta[57]),
    .outb(pe2netb[57])
  );


  cgra0_pe
  #(
    .PE_ID(59)
  )
  pe_59
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[58]),
    .branch_in(net_branch2peb[58]),
    .branch_out(pe2net_branch[58]),
    .ina(net2pea[58]),
    .inb(net2peb[58]),
    .outa(pe2neta[58]),
    .outb(pe2netb[58])
  );


  cgra0_pe
  #(
    .PE_ID(60)
  )
  pe_60
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[59]),
    .branch_in(net_branch2peb[59]),
    .branch_out(pe2net_branch[59]),
    .ina(net2pea[59]),
    .inb(net2peb[59]),
    .outa(pe2neta[59]),
    .outb(pe2netb[59])
  );


  cgra0_pe
  #(
    .PE_ID(61)
  )
  pe_61
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[60]),
    .branch_in(net_branch2peb[60]),
    .branch_out(pe2net_branch[60]),
    .ina(net2pea[60]),
    .inb(net2peb[60]),
    .outa(pe2neta[60]),
    .outb(pe2netb[60])
  );


  cgra0_pe
  #(
    .PE_ID(62)
  )
  pe_62
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[61]),
    .branch_in(net_branch2peb[61]),
    .branch_out(pe2net_branch[61]),
    .ina(net2pea[61]),
    .inb(net2peb[61]),
    .outa(pe2neta[61]),
    .outb(pe2netb[61])
  );


  cgra0_pe
  #(
    .PE_ID(63)
  )
  pe_63
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[62]),
    .branch_in(net_branch2peb[62]),
    .branch_out(pe2net_branch[62]),
    .ina(net2pea[62]),
    .inb(net2peb[62]),
    .outa(pe2neta[62]),
    .outb(pe2netb[62])
  );


  cgra0_pe
  #(
    .PE_ID(64)
  )
  pe_64
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[63]),
    .branch_in(net_branch2peb[63]),
    .branch_out(pe2net_branch[63]),
    .ina(net2pea[63]),
    .inb(net2peb[63]),
    .outa(pe2neta[63]),
    .outb(pe2netb[63])
  );


  cgra0_pe
  #(
    .PE_ID(65)
  )
  pe_65
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[64]),
    .branch_in(net_branch2peb[64]),
    .branch_out(pe2net_branch[64]),
    .ina(net2pea[64]),
    .inb(net2peb[64]),
    .outa(pe2neta[64]),
    .outb(pe2netb[64])
  );


  cgra0_pe
  #(
    .PE_ID(66)
  )
  pe_66
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[65]),
    .branch_in(net_branch2peb[65]),
    .branch_out(pe2net_branch[65]),
    .ina(net2pea[65]),
    .inb(net2peb[65]),
    .outa(pe2neta[65]),
    .outb(pe2netb[65])
  );


  cgra0_pe
  #(
    .PE_ID(67)
  )
  pe_67
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[66]),
    .branch_in(net_branch2peb[66]),
    .branch_out(pe2net_branch[66]),
    .ina(net2pea[66]),
    .inb(net2peb[66]),
    .outa(pe2neta[66]),
    .outb(pe2netb[66])
  );


  cgra0_pe
  #(
    .PE_ID(68)
  )
  pe_68
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[67]),
    .branch_in(net_branch2peb[67]),
    .branch_out(pe2net_branch[67]),
    .ina(net2pea[67]),
    .inb(net2peb[67]),
    .outa(pe2neta[67]),
    .outb(pe2netb[67])
  );


  cgra0_pe
  #(
    .PE_ID(69)
  )
  pe_69
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[68]),
    .branch_in(net_branch2peb[68]),
    .branch_out(pe2net_branch[68]),
    .ina(net2pea[68]),
    .inb(net2peb[68]),
    .outa(pe2neta[68]),
    .outb(pe2netb[68])
  );


  cgra0_pe
  #(
    .PE_ID(70)
  )
  pe_70
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[69]),
    .branch_in(net_branch2peb[69]),
    .branch_out(pe2net_branch[69]),
    .ina(net2pea[69]),
    .inb(net2peb[69]),
    .outa(pe2neta[69]),
    .outb(pe2netb[69])
  );


  cgra0_pe
  #(
    .PE_ID(71)
  )
  pe_71
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[70]),
    .branch_in(net_branch2peb[70]),
    .branch_out(pe2net_branch[70]),
    .ina(net2pea[70]),
    .inb(net2peb[70]),
    .outa(pe2neta[70]),
    .outb(pe2netb[70])
  );


  cgra0_pe
  #(
    .PE_ID(72)
  )
  pe_72
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[71]),
    .branch_in(net_branch2peb[71]),
    .branch_out(pe2net_branch[71]),
    .ina(net2pea[71]),
    .inb(net2peb[71]),
    .outa(pe2neta[71]),
    .outb(pe2netb[71])
  );


  cgra0_pe
  #(
    .PE_ID(73)
  )
  pe_73
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[72]),
    .branch_in(net_branch2peb[72]),
    .branch_out(pe2net_branch[72]),
    .ina(net2pea[72]),
    .inb(net2peb[72]),
    .outa(pe2neta[72]),
    .outb(pe2netb[72])
  );


  cgra0_pe
  #(
    .PE_ID(74)
  )
  pe_74
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[73]),
    .branch_in(net_branch2peb[73]),
    .branch_out(pe2net_branch[73]),
    .ina(net2pea[73]),
    .inb(net2peb[73]),
    .outa(pe2neta[73]),
    .outb(pe2netb[73])
  );


  cgra0_pe
  #(
    .PE_ID(75)
  )
  pe_75
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[74]),
    .branch_in(net_branch2peb[74]),
    .branch_out(pe2net_branch[74]),
    .ina(net2pea[74]),
    .inb(net2peb[74]),
    .outa(pe2neta[74]),
    .outb(pe2netb[74])
  );


  cgra0_pe
  #(
    .PE_ID(76)
  )
  pe_76
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[75]),
    .branch_in(net_branch2peb[75]),
    .branch_out(pe2net_branch[75]),
    .ina(net2pea[75]),
    .inb(net2peb[75]),
    .outa(pe2neta[75]),
    .outb(pe2netb[75])
  );


  cgra0_pe
  #(
    .PE_ID(77)
  )
  pe_77
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[76]),
    .branch_in(net_branch2peb[76]),
    .branch_out(pe2net_branch[76]),
    .ina(net2pea[76]),
    .inb(net2peb[76]),
    .outa(pe2neta[76]),
    .outb(pe2netb[76])
  );


  cgra0_pe
  #(
    .PE_ID(78)
  )
  pe_78
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[77]),
    .branch_in(net_branch2peb[77]),
    .branch_out(pe2net_branch[77]),
    .ina(net2pea[77]),
    .inb(net2peb[77]),
    .outa(pe2neta[77]),
    .outb(pe2netb[77])
  );


  cgra0_pe
  #(
    .PE_ID(79)
  )
  pe_79
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[78]),
    .branch_in(net_branch2peb[78]),
    .branch_out(pe2net_branch[78]),
    .ina(net2pea[78]),
    .inb(net2peb[78]),
    .outa(pe2neta[78]),
    .outb(pe2netb[78])
  );


  cgra0_pe
  #(
    .PE_ID(80)
  )
  pe_80
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[79]),
    .branch_in(net_branch2peb[79]),
    .branch_out(pe2net_branch[79]),
    .ina(net2pea[79]),
    .inb(net2peb[79]),
    .outa(pe2neta[79]),
    .outb(pe2netb[79])
  );


  cgra0_pe
  #(
    .PE_ID(81)
  )
  pe_81
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[80]),
    .branch_in(net_branch2peb[80]),
    .branch_out(pe2net_branch[80]),
    .ina(net2pea[80]),
    .inb(net2peb[80]),
    .outa(pe2neta[80]),
    .outb(pe2netb[80])
  );


  cgra0_pe
  #(
    .PE_ID(82)
  )
  pe_82
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[81]),
    .branch_in(net_branch2peb[81]),
    .branch_out(pe2net_branch[81]),
    .ina(net2pea[81]),
    .inb(net2peb[81]),
    .outa(pe2neta[81]),
    .outb(pe2netb[81])
  );


  cgra0_pe
  #(
    .PE_ID(83)
  )
  pe_83
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[82]),
    .branch_in(net_branch2peb[82]),
    .branch_out(pe2net_branch[82]),
    .ina(net2pea[82]),
    .inb(net2peb[82]),
    .outa(pe2neta[82]),
    .outb(pe2netb[82])
  );


  cgra0_pe
  #(
    .PE_ID(84)
  )
  pe_84
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[83]),
    .branch_in(net_branch2peb[83]),
    .branch_out(pe2net_branch[83]),
    .ina(net2pea[83]),
    .inb(net2peb[83]),
    .outa(pe2neta[83]),
    .outb(pe2netb[83])
  );


  cgra0_pe
  #(
    .PE_ID(85)
  )
  pe_85
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[84]),
    .branch_in(net_branch2peb[84]),
    .branch_out(pe2net_branch[84]),
    .ina(net2pea[84]),
    .inb(net2peb[84]),
    .outa(pe2neta[84]),
    .outb(pe2netb[84])
  );


  cgra0_pe
  #(
    .PE_ID(86)
  )
  pe_86
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[85]),
    .branch_in(net_branch2peb[85]),
    .branch_out(pe2net_branch[85]),
    .ina(net2pea[85]),
    .inb(net2peb[85]),
    .outa(pe2neta[85]),
    .outb(pe2netb[85])
  );


  cgra0_pe
  #(
    .PE_ID(87)
  )
  pe_87
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[86]),
    .branch_in(net_branch2peb[86]),
    .branch_out(pe2net_branch[86]),
    .ina(net2pea[86]),
    .inb(net2peb[86]),
    .outa(pe2neta[86]),
    .outb(pe2netb[86])
  );


  cgra0_pe
  #(
    .PE_ID(88)
  )
  pe_88
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[87]),
    .branch_in(net_branch2peb[87]),
    .branch_out(pe2net_branch[87]),
    .ina(net2pea[87]),
    .inb(net2peb[87]),
    .outa(pe2neta[87]),
    .outb(pe2netb[87])
  );


  cgra0_pe
  #(
    .PE_ID(89)
  )
  pe_89
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[88]),
    .branch_in(net_branch2peb[88]),
    .branch_out(pe2net_branch[88]),
    .ina(net2pea[88]),
    .inb(net2peb[88]),
    .outa(pe2neta[88]),
    .outb(pe2netb[88])
  );


  cgra0_pe
  #(
    .PE_ID(90)
  )
  pe_90
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[89]),
    .branch_in(net_branch2peb[89]),
    .branch_out(pe2net_branch[89]),
    .ina(net2pea[89]),
    .inb(net2peb[89]),
    .outa(pe2neta[89]),
    .outb(pe2netb[89])
  );


  cgra0_pe
  #(
    .PE_ID(91)
  )
  pe_91
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[90]),
    .branch_in(net_branch2peb[90]),
    .branch_out(pe2net_branch[90]),
    .ina(net2pea[90]),
    .inb(net2peb[90]),
    .outa(pe2neta[90]),
    .outb(pe2netb[90])
  );


  cgra0_pe
  #(
    .PE_ID(92)
  )
  pe_92
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[91]),
    .branch_in(net_branch2peb[91]),
    .branch_out(pe2net_branch[91]),
    .ina(net2pea[91]),
    .inb(net2peb[91]),
    .outa(pe2neta[91]),
    .outb(pe2netb[91])
  );


  cgra0_pe
  #(
    .PE_ID(93)
  )
  pe_93
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[92]),
    .branch_in(net_branch2peb[92]),
    .branch_out(pe2net_branch[92]),
    .ina(net2pea[92]),
    .inb(net2peb[92]),
    .outa(pe2neta[92]),
    .outb(pe2netb[92])
  );


  cgra0_pe
  #(
    .PE_ID(94)
  )
  pe_94
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[93]),
    .branch_in(net_branch2peb[93]),
    .branch_out(pe2net_branch[93]),
    .ina(net2pea[93]),
    .inb(net2peb[93]),
    .outa(pe2neta[93]),
    .outb(pe2netb[93])
  );


  cgra0_pe
  #(
    .PE_ID(95)
  )
  pe_95
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[94]),
    .branch_in(net_branch2peb[94]),
    .branch_out(pe2net_branch[94]),
    .ina(net2pea[94]),
    .inb(net2peb[94]),
    .outa(pe2neta[94]),
    .outb(pe2netb[94])
  );


  cgra0_pe
  #(
    .PE_ID(96)
  )
  pe_96
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[95]),
    .branch_in(net_branch2peb[95]),
    .branch_out(pe2net_branch[95]),
    .ina(net2pea[95]),
    .inb(net2peb[95]),
    .outa(pe2neta[95]),
    .outb(pe2netb[95])
  );


  cgra0_pe
  #(
    .PE_ID(97)
  )
  pe_97
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[96]),
    .branch_in(net_branch2peb[96]),
    .branch_out(pe2net_branch[96]),
    .ina(net2pea[96]),
    .inb(net2peb[96]),
    .outa(pe2neta[96]),
    .outb(pe2netb[96])
  );


  cgra0_pe
  #(
    .PE_ID(98)
  )
  pe_98
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[97]),
    .branch_in(net_branch2peb[97]),
    .branch_out(pe2net_branch[97]),
    .ina(net2pea[97]),
    .inb(net2peb[97]),
    .outa(pe2neta[97]),
    .outb(pe2netb[97])
  );


  cgra0_pe
  #(
    .PE_ID(99)
  )
  pe_99
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[98]),
    .branch_in(net_branch2peb[98]),
    .branch_out(pe2net_branch[98]),
    .ina(net2pea[98]),
    .inb(net2peb[98]),
    .outa(pe2neta[98]),
    .outb(pe2netb[98])
  );


  cgra0_pe
  #(
    .PE_ID(100)
  )
  pe_100
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[99]),
    .branch_in(net_branch2peb[99]),
    .branch_out(pe2net_branch[99]),
    .ina(net2pea[99]),
    .inb(net2peb[99]),
    .outa(pe2neta[99]),
    .outb(pe2netb[99])
  );


  cgra0_pe
  #(
    .PE_ID(101)
  )
  pe_101
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[100]),
    .branch_in(net_branch2peb[100]),
    .branch_out(pe2net_branch[100]),
    .ina(net2pea[100]),
    .inb(net2peb[100]),
    .outa(pe2neta[100]),
    .outb(pe2netb[100])
  );


  cgra0_pe
  #(
    .PE_ID(102)
  )
  pe_102
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[101]),
    .branch_in(net_branch2peb[101]),
    .branch_out(pe2net_branch[101]),
    .ina(net2pea[101]),
    .inb(net2peb[101]),
    .outa(pe2neta[101]),
    .outb(pe2netb[101])
  );


  cgra0_pe
  #(
    .PE_ID(103)
  )
  pe_103
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[102]),
    .branch_in(net_branch2peb[102]),
    .branch_out(pe2net_branch[102]),
    .ina(net2pea[102]),
    .inb(net2peb[102]),
    .outa(pe2neta[102]),
    .outb(pe2netb[102])
  );


  cgra0_pe
  #(
    .PE_ID(104)
  )
  pe_104
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[103]),
    .branch_in(net_branch2peb[103]),
    .branch_out(pe2net_branch[103]),
    .ina(net2pea[103]),
    .inb(net2peb[103]),
    .outa(pe2neta[103]),
    .outb(pe2netb[103])
  );


  cgra0_pe
  #(
    .PE_ID(105)
  )
  pe_105
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[104]),
    .branch_in(net_branch2peb[104]),
    .branch_out(pe2net_branch[104]),
    .ina(net2pea[104]),
    .inb(net2peb[104]),
    .outa(pe2neta[104]),
    .outb(pe2netb[104])
  );


  cgra0_pe
  #(
    .PE_ID(106)
  )
  pe_106
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[105]),
    .branch_in(net_branch2peb[105]),
    .branch_out(pe2net_branch[105]),
    .ina(net2pea[105]),
    .inb(net2peb[105]),
    .outa(pe2neta[105]),
    .outb(pe2netb[105])
  );


  cgra0_pe
  #(
    .PE_ID(107)
  )
  pe_107
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[106]),
    .branch_in(net_branch2peb[106]),
    .branch_out(pe2net_branch[106]),
    .ina(net2pea[106]),
    .inb(net2peb[106]),
    .outa(pe2neta[106]),
    .outb(pe2netb[106])
  );


  cgra0_pe
  #(
    .PE_ID(108)
  )
  pe_108
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[107]),
    .branch_in(net_branch2peb[107]),
    .branch_out(pe2net_branch[107]),
    .ina(net2pea[107]),
    .inb(net2peb[107]),
    .outa(pe2neta[107]),
    .outb(pe2netb[107])
  );


  cgra0_pe
  #(
    .PE_ID(109)
  )
  pe_109
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[108]),
    .branch_in(net_branch2peb[108]),
    .branch_out(pe2net_branch[108]),
    .ina(net2pea[108]),
    .inb(net2peb[108]),
    .outa(pe2neta[108]),
    .outb(pe2netb[108])
  );


  cgra0_pe
  #(
    .PE_ID(110)
  )
  pe_110
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[109]),
    .branch_in(net_branch2peb[109]),
    .branch_out(pe2net_branch[109]),
    .ina(net2pea[109]),
    .inb(net2peb[109]),
    .outa(pe2neta[109]),
    .outb(pe2netb[109])
  );


  cgra0_pe
  #(
    .PE_ID(111)
  )
  pe_111
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[110]),
    .branch_in(net_branch2peb[110]),
    .branch_out(pe2net_branch[110]),
    .ina(net2pea[110]),
    .inb(net2peb[110]),
    .outa(pe2neta[110]),
    .outb(pe2netb[110])
  );


  cgra0_pe
  #(
    .PE_ID(112)
  )
  pe_112
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[111]),
    .branch_in(net_branch2peb[111]),
    .branch_out(pe2net_branch[111]),
    .ina(net2pea[111]),
    .inb(net2peb[111]),
    .outa(pe2neta[111]),
    .outb(pe2netb[111])
  );


  cgra0_pe
  #(
    .PE_ID(113)
  )
  pe_113
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[112]),
    .branch_in(net_branch2peb[112]),
    .branch_out(pe2net_branch[112]),
    .ina(net2pea[112]),
    .inb(net2peb[112]),
    .outa(pe2neta[112]),
    .outb(pe2netb[112])
  );


  cgra0_pe
  #(
    .PE_ID(114)
  )
  pe_114
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[113]),
    .branch_in(net_branch2peb[113]),
    .branch_out(pe2net_branch[113]),
    .ina(net2pea[113]),
    .inb(net2peb[113]),
    .outa(pe2neta[113]),
    .outb(pe2netb[113])
  );


  cgra0_pe
  #(
    .PE_ID(115)
  )
  pe_115
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[114]),
    .branch_in(net_branch2peb[114]),
    .branch_out(pe2net_branch[114]),
    .ina(net2pea[114]),
    .inb(net2peb[114]),
    .outa(pe2neta[114]),
    .outb(pe2netb[114])
  );


  cgra0_pe
  #(
    .PE_ID(116)
  )
  pe_116
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[115]),
    .branch_in(net_branch2peb[115]),
    .branch_out(pe2net_branch[115]),
    .ina(net2pea[115]),
    .inb(net2peb[115]),
    .outa(pe2neta[115]),
    .outb(pe2netb[115])
  );


  cgra0_pe
  #(
    .PE_ID(117)
  )
  pe_117
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[116]),
    .branch_in(net_branch2peb[116]),
    .branch_out(pe2net_branch[116]),
    .ina(net2pea[116]),
    .inb(net2peb[116]),
    .outa(pe2neta[116]),
    .outb(pe2netb[116])
  );


  cgra0_pe
  #(
    .PE_ID(118)
  )
  pe_118
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[117]),
    .branch_in(net_branch2peb[117]),
    .branch_out(pe2net_branch[117]),
    .ina(net2pea[117]),
    .inb(net2peb[117]),
    .outa(pe2neta[117]),
    .outb(pe2netb[117])
  );


  cgra0_pe
  #(
    .PE_ID(119)
  )
  pe_119
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[118]),
    .branch_in(net_branch2peb[118]),
    .branch_out(pe2net_branch[118]),
    .ina(net2pea[118]),
    .inb(net2peb[118]),
    .outa(pe2neta[118]),
    .outb(pe2netb[118])
  );


  cgra0_pe
  #(
    .PE_ID(120)
  )
  pe_120
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[119]),
    .branch_in(net_branch2peb[119]),
    .branch_out(pe2net_branch[119]),
    .ina(net2pea[119]),
    .inb(net2peb[119]),
    .outa(pe2neta[119]),
    .outb(pe2netb[119])
  );


  cgra0_pe_out
  #(
    .PE_ID(121)
  )
  pe_io_out_121
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[120]),
    .branch_in(net_branch2peb[120]),
    .branch_out(pe2net_branch[120]),
    .fifo_we(fifo_out_we[0]),
    .fifo_data(fifo_out_data[15:0]),
    .ina(net2pea[120]),
    .inb(net2peb[120]),
    .outa(pe2neta[120]),
    .outb(pe2netb[120])
  );


  cgra0_pe_out
  #(
    .PE_ID(122)
  )
  pe_io_out_122
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[121]),
    .branch_in(net_branch2peb[121]),
    .branch_out(pe2net_branch[121]),
    .fifo_we(fifo_out_we[1]),
    .fifo_data(fifo_out_data[31:16]),
    .ina(net2pea[121]),
    .inb(net2peb[121]),
    .outa(pe2neta[121]),
    .outb(pe2netb[121])
  );


  cgra0_pe_out
  #(
    .PE_ID(123)
  )
  pe_io_out_123
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[122]),
    .branch_in(net_branch2peb[122]),
    .branch_out(pe2net_branch[122]),
    .fifo_we(fifo_out_we[2]),
    .fifo_data(fifo_out_data[47:32]),
    .ina(net2pea[122]),
    .inb(net2peb[122]),
    .outa(pe2neta[122]),
    .outb(pe2netb[122])
  );


  cgra0_pe_out
  #(
    .PE_ID(124)
  )
  pe_io_out_124
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[123]),
    .branch_in(net_branch2peb[123]),
    .branch_out(pe2net_branch[123]),
    .fifo_we(fifo_out_we[3]),
    .fifo_data(fifo_out_data[63:48]),
    .ina(net2pea[123]),
    .inb(net2peb[123]),
    .outa(pe2neta[123]),
    .outb(pe2netb[123])
  );


  cgra0_pe_out
  #(
    .PE_ID(125)
  )
  pe_io_out_125
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[124]),
    .branch_in(net_branch2peb[124]),
    .branch_out(pe2net_branch[124]),
    .fifo_we(fifo_out_we[4]),
    .fifo_data(fifo_out_data[79:64]),
    .ina(net2pea[124]),
    .inb(net2peb[124]),
    .outa(pe2neta[124]),
    .outb(pe2netb[124])
  );


  cgra0_pe_out
  #(
    .PE_ID(126)
  )
  pe_io_out_126
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[125]),
    .branch_in(net_branch2peb[125]),
    .branch_out(pe2net_branch[125]),
    .fifo_we(fifo_out_we[5]),
    .fifo_data(fifo_out_data[95:80]),
    .ina(net2pea[125]),
    .inb(net2peb[125]),
    .outa(pe2neta[125]),
    .outb(pe2netb[125])
  );


  cgra0_pe_out
  #(
    .PE_ID(127)
  )
  pe_io_out_127
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[126]),
    .branch_in(net_branch2peb[126]),
    .branch_out(pe2net_branch[126]),
    .fifo_we(fifo_out_we[6]),
    .fifo_data(fifo_out_data[111:96]),
    .ina(net2pea[126]),
    .inb(net2peb[126]),
    .outa(pe2neta[126]),
    .outb(pe2netb[126])
  );


  cgra0_pe_out
  #(
    .PE_ID(128)
  )
  pe_io_out_128
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .conf_bus_in(conf_bus[127]),
    .branch_in(net_branch2peb[127]),
    .branch_out(pe2net_branch[127]),
    .fifo_we(fifo_out_we[7]),
    .fifo_data(fifo_out_data[127:112]),
    .ina(net2pea[127]),
    .inb(net2peb[127]),
    .outa(pe2neta[127]),
    .outb(pe2netb[127])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_0
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[0]),
    .out(conf_bus[1])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_1
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[1]),
    .out(conf_bus[2])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_2
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[2]),
    .out(conf_bus[3])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_3
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[3]),
    .out(conf_bus[4])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_4
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[4]),
    .out(conf_bus[5])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_5
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[5]),
    .out(conf_bus[6])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_6
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[6]),
    .out(conf_bus[7])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_7
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[7]),
    .out(conf_bus[8])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_8
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[8]),
    .out(conf_bus[9])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_9
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[9]),
    .out(conf_bus[10])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_10
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[10]),
    .out(conf_bus[11])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_11
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[11]),
    .out(conf_bus[12])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_12
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[12]),
    .out(conf_bus[13])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_13
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[13]),
    .out(conf_bus[14])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_14
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[14]),
    .out(conf_bus[15])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_15
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[15]),
    .out(conf_bus[16])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_16
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[16]),
    .out(conf_bus[17])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_17
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[17]),
    .out(conf_bus[18])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_18
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[18]),
    .out(conf_bus[19])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_19
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[19]),
    .out(conf_bus[20])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_20
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[20]),
    .out(conf_bus[21])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_21
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[21]),
    .out(conf_bus[22])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_22
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[22]),
    .out(conf_bus[23])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_23
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[23]),
    .out(conf_bus[24])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_24
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[24]),
    .out(conf_bus[25])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_25
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[25]),
    .out(conf_bus[26])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_26
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[26]),
    .out(conf_bus[27])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_27
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[27]),
    .out(conf_bus[28])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_28
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[28]),
    .out(conf_bus[29])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_29
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[29]),
    .out(conf_bus[30])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_30
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[30]),
    .out(conf_bus[31])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_31
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[31]),
    .out(conf_bus[32])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_32
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[32]),
    .out(conf_bus[33])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_33
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[33]),
    .out(conf_bus[34])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_34
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[34]),
    .out(conf_bus[35])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_35
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[35]),
    .out(conf_bus[36])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_36
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[36]),
    .out(conf_bus[37])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_37
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[37]),
    .out(conf_bus[38])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_38
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[38]),
    .out(conf_bus[39])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_39
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[39]),
    .out(conf_bus[40])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_40
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[40]),
    .out(conf_bus[41])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_41
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[41]),
    .out(conf_bus[42])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_42
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[42]),
    .out(conf_bus[43])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_43
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[43]),
    .out(conf_bus[44])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_44
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[44]),
    .out(conf_bus[45])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_45
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[45]),
    .out(conf_bus[46])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_46
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[46]),
    .out(conf_bus[47])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_47
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[47]),
    .out(conf_bus[48])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_48
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[48]),
    .out(conf_bus[49])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_49
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[49]),
    .out(conf_bus[50])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_50
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[50]),
    .out(conf_bus[51])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_51
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[51]),
    .out(conf_bus[52])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_52
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[52]),
    .out(conf_bus[53])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_53
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[53]),
    .out(conf_bus[54])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_54
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[54]),
    .out(conf_bus[55])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_55
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[55]),
    .out(conf_bus[56])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_56
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[56]),
    .out(conf_bus[57])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_57
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[57]),
    .out(conf_bus[58])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_58
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[58]),
    .out(conf_bus[59])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_59
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[59]),
    .out(conf_bus[60])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_60
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[60]),
    .out(conf_bus[61])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_61
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[61]),
    .out(conf_bus[62])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_62
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[62]),
    .out(conf_bus[63])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_63
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[63]),
    .out(conf_bus[64])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_64
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[64]),
    .out(conf_bus[65])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_65
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[65]),
    .out(conf_bus[66])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_66
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[66]),
    .out(conf_bus[67])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_67
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[67]),
    .out(conf_bus[68])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_68
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[68]),
    .out(conf_bus[69])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_69
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[69]),
    .out(conf_bus[70])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_70
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[70]),
    .out(conf_bus[71])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_71
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[71]),
    .out(conf_bus[72])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_72
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[72]),
    .out(conf_bus[73])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_73
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[73]),
    .out(conf_bus[74])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_74
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[74]),
    .out(conf_bus[75])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_75
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[75]),
    .out(conf_bus[76])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_76
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[76]),
    .out(conf_bus[77])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_77
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[77]),
    .out(conf_bus[78])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_78
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[78]),
    .out(conf_bus[79])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_79
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[79]),
    .out(conf_bus[80])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_80
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[80]),
    .out(conf_bus[81])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_81
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[81]),
    .out(conf_bus[82])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_82
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[82]),
    .out(conf_bus[83])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_83
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[83]),
    .out(conf_bus[84])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_84
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[84]),
    .out(conf_bus[85])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_85
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[85]),
    .out(conf_bus[86])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_86
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[86]),
    .out(conf_bus[87])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_87
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[87]),
    .out(conf_bus[88])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_88
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[88]),
    .out(conf_bus[89])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_89
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[89]),
    .out(conf_bus[90])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_90
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[90]),
    .out(conf_bus[91])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_91
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[91]),
    .out(conf_bus[92])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_92
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[92]),
    .out(conf_bus[93])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_93
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[93]),
    .out(conf_bus[94])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_94
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[94]),
    .out(conf_bus[95])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_95
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[95]),
    .out(conf_bus[96])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_96
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[96]),
    .out(conf_bus[97])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_97
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[97]),
    .out(conf_bus[98])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_98
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[98]),
    .out(conf_bus[99])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_99
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[99]),
    .out(conf_bus[100])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_100
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[100]),
    .out(conf_bus[101])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_101
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[101]),
    .out(conf_bus[102])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_102
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[102]),
    .out(conf_bus[103])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_103
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[103]),
    .out(conf_bus[104])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_104
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[104]),
    .out(conf_bus[105])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_105
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[105]),
    .out(conf_bus[106])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_106
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[106]),
    .out(conf_bus[107])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_107
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[107]),
    .out(conf_bus[108])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_108
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[108]),
    .out(conf_bus[109])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_109
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[109]),
    .out(conf_bus[110])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_110
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[110]),
    .out(conf_bus[111])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_111
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[111]),
    .out(conf_bus[112])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_112
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[112]),
    .out(conf_bus[113])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_113
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[113]),
    .out(conf_bus[114])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_114
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[114]),
    .out(conf_bus[115])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_115
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[115]),
    .out(conf_bus[116])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_116
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[116]),
    .out(conf_bus[117])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_117
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[117]),
    .out(conf_bus[118])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_118
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[118]),
    .out(conf_bus[119])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_119
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[119]),
    .out(conf_bus[120])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_120
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[120]),
    .out(conf_bus[121])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_121
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[121]),
    .out(conf_bus[122])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_122
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[122]),
    .out(conf_bus[123])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_123
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[123]),
    .out(conf_bus[124])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_124
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[124]),
    .out(conf_bus[125])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_125
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[125]),
    .out(conf_bus[126])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_126
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[126]),
    .out(conf_bus[127])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  conf_bus_reg_127
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(conf_bus[127]),
    .out(conf_bus[128])
  );


  omega256x256_8_1_1
  #(
    .WIDTH(16),
    .PIPE_EXTRA(0)
  )
  net
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .net_conf_bus_in(conf_bus[128]),
    .in0(pe2neta[0]),
    .in1(pe2netb[0]),
    .in2(pe2neta[1]),
    .in3(pe2netb[1]),
    .in4(pe2neta[2]),
    .in5(pe2netb[2]),
    .in6(pe2neta[3]),
    .in7(pe2netb[3]),
    .in8(pe2neta[4]),
    .in9(pe2netb[4]),
    .in10(pe2neta[5]),
    .in11(pe2netb[5]),
    .in12(pe2neta[6]),
    .in13(pe2netb[6]),
    .in14(pe2neta[7]),
    .in15(pe2netb[7]),
    .in16(pe2neta[8]),
    .in17(pe2netb[8]),
    .in18(pe2neta[9]),
    .in19(pe2netb[9]),
    .in20(pe2neta[10]),
    .in21(pe2netb[10]),
    .in22(pe2neta[11]),
    .in23(pe2netb[11]),
    .in24(pe2neta[12]),
    .in25(pe2netb[12]),
    .in26(pe2neta[13]),
    .in27(pe2netb[13]),
    .in28(pe2neta[14]),
    .in29(pe2netb[14]),
    .in30(pe2neta[15]),
    .in31(pe2netb[15]),
    .in32(pe2neta[16]),
    .in33(pe2netb[16]),
    .in34(pe2neta[17]),
    .in35(pe2netb[17]),
    .in36(pe2neta[18]),
    .in37(pe2netb[18]),
    .in38(pe2neta[19]),
    .in39(pe2netb[19]),
    .in40(pe2neta[20]),
    .in41(pe2netb[20]),
    .in42(pe2neta[21]),
    .in43(pe2netb[21]),
    .in44(pe2neta[22]),
    .in45(pe2netb[22]),
    .in46(pe2neta[23]),
    .in47(pe2netb[23]),
    .in48(pe2neta[24]),
    .in49(pe2netb[24]),
    .in50(pe2neta[25]),
    .in51(pe2netb[25]),
    .in52(pe2neta[26]),
    .in53(pe2netb[26]),
    .in54(pe2neta[27]),
    .in55(pe2netb[27]),
    .in56(pe2neta[28]),
    .in57(pe2netb[28]),
    .in58(pe2neta[29]),
    .in59(pe2netb[29]),
    .in60(pe2neta[30]),
    .in61(pe2netb[30]),
    .in62(pe2neta[31]),
    .in63(pe2netb[31]),
    .in64(pe2neta[32]),
    .in65(pe2netb[32]),
    .in66(pe2neta[33]),
    .in67(pe2netb[33]),
    .in68(pe2neta[34]),
    .in69(pe2netb[34]),
    .in70(pe2neta[35]),
    .in71(pe2netb[35]),
    .in72(pe2neta[36]),
    .in73(pe2netb[36]),
    .in74(pe2neta[37]),
    .in75(pe2netb[37]),
    .in76(pe2neta[38]),
    .in77(pe2netb[38]),
    .in78(pe2neta[39]),
    .in79(pe2netb[39]),
    .in80(pe2neta[40]),
    .in81(pe2netb[40]),
    .in82(pe2neta[41]),
    .in83(pe2netb[41]),
    .in84(pe2neta[42]),
    .in85(pe2netb[42]),
    .in86(pe2neta[43]),
    .in87(pe2netb[43]),
    .in88(pe2neta[44]),
    .in89(pe2netb[44]),
    .in90(pe2neta[45]),
    .in91(pe2netb[45]),
    .in92(pe2neta[46]),
    .in93(pe2netb[46]),
    .in94(pe2neta[47]),
    .in95(pe2netb[47]),
    .in96(pe2neta[48]),
    .in97(pe2netb[48]),
    .in98(pe2neta[49]),
    .in99(pe2netb[49]),
    .in100(pe2neta[50]),
    .in101(pe2netb[50]),
    .in102(pe2neta[51]),
    .in103(pe2netb[51]),
    .in104(pe2neta[52]),
    .in105(pe2netb[52]),
    .in106(pe2neta[53]),
    .in107(pe2netb[53]),
    .in108(pe2neta[54]),
    .in109(pe2netb[54]),
    .in110(pe2neta[55]),
    .in111(pe2netb[55]),
    .in112(pe2neta[56]),
    .in113(pe2netb[56]),
    .in114(pe2neta[57]),
    .in115(pe2netb[57]),
    .in116(pe2neta[58]),
    .in117(pe2netb[58]),
    .in118(pe2neta[59]),
    .in119(pe2netb[59]),
    .in120(pe2neta[60]),
    .in121(pe2netb[60]),
    .in122(pe2neta[61]),
    .in123(pe2netb[61]),
    .in124(pe2neta[62]),
    .in125(pe2netb[62]),
    .in126(pe2neta[63]),
    .in127(pe2netb[63]),
    .in128(pe2neta[64]),
    .in129(pe2netb[64]),
    .in130(pe2neta[65]),
    .in131(pe2netb[65]),
    .in132(pe2neta[66]),
    .in133(pe2netb[66]),
    .in134(pe2neta[67]),
    .in135(pe2netb[67]),
    .in136(pe2neta[68]),
    .in137(pe2netb[68]),
    .in138(pe2neta[69]),
    .in139(pe2netb[69]),
    .in140(pe2neta[70]),
    .in141(pe2netb[70]),
    .in142(pe2neta[71]),
    .in143(pe2netb[71]),
    .in144(pe2neta[72]),
    .in145(pe2netb[72]),
    .in146(pe2neta[73]),
    .in147(pe2netb[73]),
    .in148(pe2neta[74]),
    .in149(pe2netb[74]),
    .in150(pe2neta[75]),
    .in151(pe2netb[75]),
    .in152(pe2neta[76]),
    .in153(pe2netb[76]),
    .in154(pe2neta[77]),
    .in155(pe2netb[77]),
    .in156(pe2neta[78]),
    .in157(pe2netb[78]),
    .in158(pe2neta[79]),
    .in159(pe2netb[79]),
    .in160(pe2neta[80]),
    .in161(pe2netb[80]),
    .in162(pe2neta[81]),
    .in163(pe2netb[81]),
    .in164(pe2neta[82]),
    .in165(pe2netb[82]),
    .in166(pe2neta[83]),
    .in167(pe2netb[83]),
    .in168(pe2neta[84]),
    .in169(pe2netb[84]),
    .in170(pe2neta[85]),
    .in171(pe2netb[85]),
    .in172(pe2neta[86]),
    .in173(pe2netb[86]),
    .in174(pe2neta[87]),
    .in175(pe2netb[87]),
    .in176(pe2neta[88]),
    .in177(pe2netb[88]),
    .in178(pe2neta[89]),
    .in179(pe2netb[89]),
    .in180(pe2neta[90]),
    .in181(pe2netb[90]),
    .in182(pe2neta[91]),
    .in183(pe2netb[91]),
    .in184(pe2neta[92]),
    .in185(pe2netb[92]),
    .in186(pe2neta[93]),
    .in187(pe2netb[93]),
    .in188(pe2neta[94]),
    .in189(pe2netb[94]),
    .in190(pe2neta[95]),
    .in191(pe2netb[95]),
    .in192(pe2neta[96]),
    .in193(pe2netb[96]),
    .in194(pe2neta[97]),
    .in195(pe2netb[97]),
    .in196(pe2neta[98]),
    .in197(pe2netb[98]),
    .in198(pe2neta[99]),
    .in199(pe2netb[99]),
    .in200(pe2neta[100]),
    .in201(pe2netb[100]),
    .in202(pe2neta[101]),
    .in203(pe2netb[101]),
    .in204(pe2neta[102]),
    .in205(pe2netb[102]),
    .in206(pe2neta[103]),
    .in207(pe2netb[103]),
    .in208(pe2neta[104]),
    .in209(pe2netb[104]),
    .in210(pe2neta[105]),
    .in211(pe2netb[105]),
    .in212(pe2neta[106]),
    .in213(pe2netb[106]),
    .in214(pe2neta[107]),
    .in215(pe2netb[107]),
    .in216(pe2neta[108]),
    .in217(pe2netb[108]),
    .in218(pe2neta[109]),
    .in219(pe2netb[109]),
    .in220(pe2neta[110]),
    .in221(pe2netb[110]),
    .in222(pe2neta[111]),
    .in223(pe2netb[111]),
    .in224(pe2neta[112]),
    .in225(pe2netb[112]),
    .in226(pe2neta[113]),
    .in227(pe2netb[113]),
    .in228(pe2neta[114]),
    .in229(pe2netb[114]),
    .in230(pe2neta[115]),
    .in231(pe2netb[115]),
    .in232(pe2neta[116]),
    .in233(pe2netb[116]),
    .in234(pe2neta[117]),
    .in235(pe2netb[117]),
    .in236(pe2neta[118]),
    .in237(pe2netb[118]),
    .in238(pe2neta[119]),
    .in239(pe2netb[119]),
    .in240(pe2neta[120]),
    .in241(pe2netb[120]),
    .in242(pe2neta[121]),
    .in243(pe2netb[121]),
    .in244(pe2neta[122]),
    .in245(pe2netb[122]),
    .in246(pe2neta[123]),
    .in247(pe2netb[123]),
    .in248(pe2neta[124]),
    .in249(pe2netb[124]),
    .in250(pe2neta[125]),
    .in251(pe2netb[125]),
    .in252(pe2neta[126]),
    .in253(pe2netb[126]),
    .in254(pe2neta[127]),
    .in255(pe2netb[127]),
    .out0(net2pea[0]),
    .out1(net2peb[0]),
    .out2(net2pea[1]),
    .out3(net2peb[1]),
    .out4(net2pea[2]),
    .out5(net2peb[2]),
    .out6(net2pea[3]),
    .out7(net2peb[3]),
    .out8(net2pea[4]),
    .out9(net2peb[4]),
    .out10(net2pea[5]),
    .out11(net2peb[5]),
    .out12(net2pea[6]),
    .out13(net2peb[6]),
    .out14(net2pea[7]),
    .out15(net2peb[7]),
    .out16(net2pea[8]),
    .out17(net2peb[8]),
    .out18(net2pea[9]),
    .out19(net2peb[9]),
    .out20(net2pea[10]),
    .out21(net2peb[10]),
    .out22(net2pea[11]),
    .out23(net2peb[11]),
    .out24(net2pea[12]),
    .out25(net2peb[12]),
    .out26(net2pea[13]),
    .out27(net2peb[13]),
    .out28(net2pea[14]),
    .out29(net2peb[14]),
    .out30(net2pea[15]),
    .out31(net2peb[15]),
    .out32(net2pea[16]),
    .out33(net2peb[16]),
    .out34(net2pea[17]),
    .out35(net2peb[17]),
    .out36(net2pea[18]),
    .out37(net2peb[18]),
    .out38(net2pea[19]),
    .out39(net2peb[19]),
    .out40(net2pea[20]),
    .out41(net2peb[20]),
    .out42(net2pea[21]),
    .out43(net2peb[21]),
    .out44(net2pea[22]),
    .out45(net2peb[22]),
    .out46(net2pea[23]),
    .out47(net2peb[23]),
    .out48(net2pea[24]),
    .out49(net2peb[24]),
    .out50(net2pea[25]),
    .out51(net2peb[25]),
    .out52(net2pea[26]),
    .out53(net2peb[26]),
    .out54(net2pea[27]),
    .out55(net2peb[27]),
    .out56(net2pea[28]),
    .out57(net2peb[28]),
    .out58(net2pea[29]),
    .out59(net2peb[29]),
    .out60(net2pea[30]),
    .out61(net2peb[30]),
    .out62(net2pea[31]),
    .out63(net2peb[31]),
    .out64(net2pea[32]),
    .out65(net2peb[32]),
    .out66(net2pea[33]),
    .out67(net2peb[33]),
    .out68(net2pea[34]),
    .out69(net2peb[34]),
    .out70(net2pea[35]),
    .out71(net2peb[35]),
    .out72(net2pea[36]),
    .out73(net2peb[36]),
    .out74(net2pea[37]),
    .out75(net2peb[37]),
    .out76(net2pea[38]),
    .out77(net2peb[38]),
    .out78(net2pea[39]),
    .out79(net2peb[39]),
    .out80(net2pea[40]),
    .out81(net2peb[40]),
    .out82(net2pea[41]),
    .out83(net2peb[41]),
    .out84(net2pea[42]),
    .out85(net2peb[42]),
    .out86(net2pea[43]),
    .out87(net2peb[43]),
    .out88(net2pea[44]),
    .out89(net2peb[44]),
    .out90(net2pea[45]),
    .out91(net2peb[45]),
    .out92(net2pea[46]),
    .out93(net2peb[46]),
    .out94(net2pea[47]),
    .out95(net2peb[47]),
    .out96(net2pea[48]),
    .out97(net2peb[48]),
    .out98(net2pea[49]),
    .out99(net2peb[49]),
    .out100(net2pea[50]),
    .out101(net2peb[50]),
    .out102(net2pea[51]),
    .out103(net2peb[51]),
    .out104(net2pea[52]),
    .out105(net2peb[52]),
    .out106(net2pea[53]),
    .out107(net2peb[53]),
    .out108(net2pea[54]),
    .out109(net2peb[54]),
    .out110(net2pea[55]),
    .out111(net2peb[55]),
    .out112(net2pea[56]),
    .out113(net2peb[56]),
    .out114(net2pea[57]),
    .out115(net2peb[57]),
    .out116(net2pea[58]),
    .out117(net2peb[58]),
    .out118(net2pea[59]),
    .out119(net2peb[59]),
    .out120(net2pea[60]),
    .out121(net2peb[60]),
    .out122(net2pea[61]),
    .out123(net2peb[61]),
    .out124(net2pea[62]),
    .out125(net2peb[62]),
    .out126(net2pea[63]),
    .out127(net2peb[63]),
    .out128(net2pea[64]),
    .out129(net2peb[64]),
    .out130(net2pea[65]),
    .out131(net2peb[65]),
    .out132(net2pea[66]),
    .out133(net2peb[66]),
    .out134(net2pea[67]),
    .out135(net2peb[67]),
    .out136(net2pea[68]),
    .out137(net2peb[68]),
    .out138(net2pea[69]),
    .out139(net2peb[69]),
    .out140(net2pea[70]),
    .out141(net2peb[70]),
    .out142(net2pea[71]),
    .out143(net2peb[71]),
    .out144(net2pea[72]),
    .out145(net2peb[72]),
    .out146(net2pea[73]),
    .out147(net2peb[73]),
    .out148(net2pea[74]),
    .out149(net2peb[74]),
    .out150(net2pea[75]),
    .out151(net2peb[75]),
    .out152(net2pea[76]),
    .out153(net2peb[76]),
    .out154(net2pea[77]),
    .out155(net2peb[77]),
    .out156(net2pea[78]),
    .out157(net2peb[78]),
    .out158(net2pea[79]),
    .out159(net2peb[79]),
    .out160(net2pea[80]),
    .out161(net2peb[80]),
    .out162(net2pea[81]),
    .out163(net2peb[81]),
    .out164(net2pea[82]),
    .out165(net2peb[82]),
    .out166(net2pea[83]),
    .out167(net2peb[83]),
    .out168(net2pea[84]),
    .out169(net2peb[84]),
    .out170(net2pea[85]),
    .out171(net2peb[85]),
    .out172(net2pea[86]),
    .out173(net2peb[86]),
    .out174(net2pea[87]),
    .out175(net2peb[87]),
    .out176(net2pea[88]),
    .out177(net2peb[88]),
    .out178(net2pea[89]),
    .out179(net2peb[89]),
    .out180(net2pea[90]),
    .out181(net2peb[90]),
    .out182(net2pea[91]),
    .out183(net2peb[91]),
    .out184(net2pea[92]),
    .out185(net2peb[92]),
    .out186(net2pea[93]),
    .out187(net2peb[93]),
    .out188(net2pea[94]),
    .out189(net2peb[94]),
    .out190(net2pea[95]),
    .out191(net2peb[95]),
    .out192(net2pea[96]),
    .out193(net2peb[96]),
    .out194(net2pea[97]),
    .out195(net2peb[97]),
    .out196(net2pea[98]),
    .out197(net2peb[98]),
    .out198(net2pea[99]),
    .out199(net2peb[99]),
    .out200(net2pea[100]),
    .out201(net2peb[100]),
    .out202(net2pea[101]),
    .out203(net2peb[101]),
    .out204(net2pea[102]),
    .out205(net2peb[102]),
    .out206(net2pea[103]),
    .out207(net2peb[103]),
    .out208(net2pea[104]),
    .out209(net2peb[104]),
    .out210(net2pea[105]),
    .out211(net2peb[105]),
    .out212(net2pea[106]),
    .out213(net2peb[106]),
    .out214(net2pea[107]),
    .out215(net2peb[107]),
    .out216(net2pea[108]),
    .out217(net2peb[108]),
    .out218(net2pea[109]),
    .out219(net2peb[109]),
    .out220(net2pea[110]),
    .out221(net2peb[110]),
    .out222(net2pea[111]),
    .out223(net2peb[111]),
    .out224(net2pea[112]),
    .out225(net2peb[112]),
    .out226(net2pea[113]),
    .out227(net2peb[113]),
    .out228(net2pea[114]),
    .out229(net2peb[114]),
    .out230(net2pea[115]),
    .out231(net2peb[115]),
    .out232(net2pea[116]),
    .out233(net2peb[116]),
    .out234(net2pea[117]),
    .out235(net2peb[117]),
    .out236(net2pea[118]),
    .out237(net2peb[118]),
    .out238(net2pea[119]),
    .out239(net2peb[119]),
    .out240(net2pea[120]),
    .out241(net2peb[120]),
    .out242(net2pea[121]),
    .out243(net2peb[121]),
    .out244(net2pea[122]),
    .out245(net2peb[122]),
    .out246(net2pea[123]),
    .out247(net2peb[123]),
    .out248(net2pea[124]),
    .out249(net2peb[124]),
    .out250(net2pea[125]),
    .out251(net2peb[125]),
    .out252(net2pea[126]),
    .out253(net2peb[126]),
    .out254(net2pea[127]),
    .out255(net2peb[127])
  );


  omega_branch128x128_8_1_1
  #(
    .WIDTH(1),
    .PIPE_EXTRA(0)
  )
  net_branch
  (
    .clk(clk),
    .rst(rst),
    .en(en),
    .net_conf_bus_in(conf_bus[128]),
    .in0(pe2net_branch[0]),
    .in1(pe2net_branch[1]),
    .in2(pe2net_branch[2]),
    .in3(pe2net_branch[3]),
    .in4(pe2net_branch[4]),
    .in5(pe2net_branch[5]),
    .in6(pe2net_branch[6]),
    .in7(pe2net_branch[7]),
    .in8(pe2net_branch[8]),
    .in9(pe2net_branch[9]),
    .in10(pe2net_branch[10]),
    .in11(pe2net_branch[11]),
    .in12(pe2net_branch[12]),
    .in13(pe2net_branch[13]),
    .in14(pe2net_branch[14]),
    .in15(pe2net_branch[15]),
    .in16(pe2net_branch[16]),
    .in17(pe2net_branch[17]),
    .in18(pe2net_branch[18]),
    .in19(pe2net_branch[19]),
    .in20(pe2net_branch[20]),
    .in21(pe2net_branch[21]),
    .in22(pe2net_branch[22]),
    .in23(pe2net_branch[23]),
    .in24(pe2net_branch[24]),
    .in25(pe2net_branch[25]),
    .in26(pe2net_branch[26]),
    .in27(pe2net_branch[27]),
    .in28(pe2net_branch[28]),
    .in29(pe2net_branch[29]),
    .in30(pe2net_branch[30]),
    .in31(pe2net_branch[31]),
    .in32(pe2net_branch[32]),
    .in33(pe2net_branch[33]),
    .in34(pe2net_branch[34]),
    .in35(pe2net_branch[35]),
    .in36(pe2net_branch[36]),
    .in37(pe2net_branch[37]),
    .in38(pe2net_branch[38]),
    .in39(pe2net_branch[39]),
    .in40(pe2net_branch[40]),
    .in41(pe2net_branch[41]),
    .in42(pe2net_branch[42]),
    .in43(pe2net_branch[43]),
    .in44(pe2net_branch[44]),
    .in45(pe2net_branch[45]),
    .in46(pe2net_branch[46]),
    .in47(pe2net_branch[47]),
    .in48(pe2net_branch[48]),
    .in49(pe2net_branch[49]),
    .in50(pe2net_branch[50]),
    .in51(pe2net_branch[51]),
    .in52(pe2net_branch[52]),
    .in53(pe2net_branch[53]),
    .in54(pe2net_branch[54]),
    .in55(pe2net_branch[55]),
    .in56(pe2net_branch[56]),
    .in57(pe2net_branch[57]),
    .in58(pe2net_branch[58]),
    .in59(pe2net_branch[59]),
    .in60(pe2net_branch[60]),
    .in61(pe2net_branch[61]),
    .in62(pe2net_branch[62]),
    .in63(pe2net_branch[63]),
    .in64(pe2net_branch[64]),
    .in65(pe2net_branch[65]),
    .in66(pe2net_branch[66]),
    .in67(pe2net_branch[67]),
    .in68(pe2net_branch[68]),
    .in69(pe2net_branch[69]),
    .in70(pe2net_branch[70]),
    .in71(pe2net_branch[71]),
    .in72(pe2net_branch[72]),
    .in73(pe2net_branch[73]),
    .in74(pe2net_branch[74]),
    .in75(pe2net_branch[75]),
    .in76(pe2net_branch[76]),
    .in77(pe2net_branch[77]),
    .in78(pe2net_branch[78]),
    .in79(pe2net_branch[79]),
    .in80(pe2net_branch[80]),
    .in81(pe2net_branch[81]),
    .in82(pe2net_branch[82]),
    .in83(pe2net_branch[83]),
    .in84(pe2net_branch[84]),
    .in85(pe2net_branch[85]),
    .in86(pe2net_branch[86]),
    .in87(pe2net_branch[87]),
    .in88(pe2net_branch[88]),
    .in89(pe2net_branch[89]),
    .in90(pe2net_branch[90]),
    .in91(pe2net_branch[91]),
    .in92(pe2net_branch[92]),
    .in93(pe2net_branch[93]),
    .in94(pe2net_branch[94]),
    .in95(pe2net_branch[95]),
    .in96(pe2net_branch[96]),
    .in97(pe2net_branch[97]),
    .in98(pe2net_branch[98]),
    .in99(pe2net_branch[99]),
    .in100(pe2net_branch[100]),
    .in101(pe2net_branch[101]),
    .in102(pe2net_branch[102]),
    .in103(pe2net_branch[103]),
    .in104(pe2net_branch[104]),
    .in105(pe2net_branch[105]),
    .in106(pe2net_branch[106]),
    .in107(pe2net_branch[107]),
    .in108(pe2net_branch[108]),
    .in109(pe2net_branch[109]),
    .in110(pe2net_branch[110]),
    .in111(pe2net_branch[111]),
    .in112(pe2net_branch[112]),
    .in113(pe2net_branch[113]),
    .in114(pe2net_branch[114]),
    .in115(pe2net_branch[115]),
    .in116(pe2net_branch[116]),
    .in117(pe2net_branch[117]),
    .in118(pe2net_branch[118]),
    .in119(pe2net_branch[119]),
    .in120(pe2net_branch[120]),
    .in121(pe2net_branch[121]),
    .in122(pe2net_branch[122]),
    .in123(pe2net_branch[123]),
    .in124(pe2net_branch[124]),
    .in125(pe2net_branch[125]),
    .in126(pe2net_branch[126]),
    .in127(pe2net_branch[127]),
    .out0(net_branch2peb[0]),
    .out1(net_branch2peb[1]),
    .out2(net_branch2peb[2]),
    .out3(net_branch2peb[3]),
    .out4(net_branch2peb[4]),
    .out5(net_branch2peb[5]),
    .out6(net_branch2peb[6]),
    .out7(net_branch2peb[7]),
    .out8(net_branch2peb[8]),
    .out9(net_branch2peb[9]),
    .out10(net_branch2peb[10]),
    .out11(net_branch2peb[11]),
    .out12(net_branch2peb[12]),
    .out13(net_branch2peb[13]),
    .out14(net_branch2peb[14]),
    .out15(net_branch2peb[15]),
    .out16(net_branch2peb[16]),
    .out17(net_branch2peb[17]),
    .out18(net_branch2peb[18]),
    .out19(net_branch2peb[19]),
    .out20(net_branch2peb[20]),
    .out21(net_branch2peb[21]),
    .out22(net_branch2peb[22]),
    .out23(net_branch2peb[23]),
    .out24(net_branch2peb[24]),
    .out25(net_branch2peb[25]),
    .out26(net_branch2peb[26]),
    .out27(net_branch2peb[27]),
    .out28(net_branch2peb[28]),
    .out29(net_branch2peb[29]),
    .out30(net_branch2peb[30]),
    .out31(net_branch2peb[31]),
    .out32(net_branch2peb[32]),
    .out33(net_branch2peb[33]),
    .out34(net_branch2peb[34]),
    .out35(net_branch2peb[35]),
    .out36(net_branch2peb[36]),
    .out37(net_branch2peb[37]),
    .out38(net_branch2peb[38]),
    .out39(net_branch2peb[39]),
    .out40(net_branch2peb[40]),
    .out41(net_branch2peb[41]),
    .out42(net_branch2peb[42]),
    .out43(net_branch2peb[43]),
    .out44(net_branch2peb[44]),
    .out45(net_branch2peb[45]),
    .out46(net_branch2peb[46]),
    .out47(net_branch2peb[47]),
    .out48(net_branch2peb[48]),
    .out49(net_branch2peb[49]),
    .out50(net_branch2peb[50]),
    .out51(net_branch2peb[51]),
    .out52(net_branch2peb[52]),
    .out53(net_branch2peb[53]),
    .out54(net_branch2peb[54]),
    .out55(net_branch2peb[55]),
    .out56(net_branch2peb[56]),
    .out57(net_branch2peb[57]),
    .out58(net_branch2peb[58]),
    .out59(net_branch2peb[59]),
    .out60(net_branch2peb[60]),
    .out61(net_branch2peb[61]),
    .out62(net_branch2peb[62]),
    .out63(net_branch2peb[63]),
    .out64(net_branch2peb[64]),
    .out65(net_branch2peb[65]),
    .out66(net_branch2peb[66]),
    .out67(net_branch2peb[67]),
    .out68(net_branch2peb[68]),
    .out69(net_branch2peb[69]),
    .out70(net_branch2peb[70]),
    .out71(net_branch2peb[71]),
    .out72(net_branch2peb[72]),
    .out73(net_branch2peb[73]),
    .out74(net_branch2peb[74]),
    .out75(net_branch2peb[75]),
    .out76(net_branch2peb[76]),
    .out77(net_branch2peb[77]),
    .out78(net_branch2peb[78]),
    .out79(net_branch2peb[79]),
    .out80(net_branch2peb[80]),
    .out81(net_branch2peb[81]),
    .out82(net_branch2peb[82]),
    .out83(net_branch2peb[83]),
    .out84(net_branch2peb[84]),
    .out85(net_branch2peb[85]),
    .out86(net_branch2peb[86]),
    .out87(net_branch2peb[87]),
    .out88(net_branch2peb[88]),
    .out89(net_branch2peb[89]),
    .out90(net_branch2peb[90]),
    .out91(net_branch2peb[91]),
    .out92(net_branch2peb[92]),
    .out93(net_branch2peb[93]),
    .out94(net_branch2peb[94]),
    .out95(net_branch2peb[95]),
    .out96(net_branch2peb[96]),
    .out97(net_branch2peb[97]),
    .out98(net_branch2peb[98]),
    .out99(net_branch2peb[99]),
    .out100(net_branch2peb[100]),
    .out101(net_branch2peb[101]),
    .out102(net_branch2peb[102]),
    .out103(net_branch2peb[103]),
    .out104(net_branch2peb[104]),
    .out105(net_branch2peb[105]),
    .out106(net_branch2peb[106]),
    .out107(net_branch2peb[107]),
    .out108(net_branch2peb[108]),
    .out109(net_branch2peb[109]),
    .out110(net_branch2peb[110]),
    .out111(net_branch2peb[111]),
    .out112(net_branch2peb[112]),
    .out113(net_branch2peb[113]),
    .out114(net_branch2peb[114]),
    .out115(net_branch2peb[115]),
    .out116(net_branch2peb[116]),
    .out117(net_branch2peb[117]),
    .out118(net_branch2peb[118]),
    .out119(net_branch2peb[119]),
    .out120(net_branch2peb[120]),
    .out121(net_branch2peb[121]),
    .out122(net_branch2peb[122]),
    .out123(net_branch2peb[123]),
    .out124(net_branch2peb[124]),
    .out125(net_branch2peb[125]),
    .out126(net_branch2peb[126]),
    .out127(net_branch2peb[127])
  );

endmodule