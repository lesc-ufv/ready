module omega_branch128x128_8_1_1 #
(
  parameter WIDTH = 16,
  parameter PIPE_EXTRA = 0
)
(
  input clk,
  input rst,
  input en,
  input [64-1:0] net_conf_bus_in,
  input [WIDTH-1:0] in0,
  input [WIDTH-1:0] in1,
  input [WIDTH-1:0] in2,
  input [WIDTH-1:0] in3,
  input [WIDTH-1:0] in4,
  input [WIDTH-1:0] in5,
  input [WIDTH-1:0] in6,
  input [WIDTH-1:0] in7,
  input [WIDTH-1:0] in8,
  input [WIDTH-1:0] in9,
  input [WIDTH-1:0] in10,
  input [WIDTH-1:0] in11,
  input [WIDTH-1:0] in12,
  input [WIDTH-1:0] in13,
  input [WIDTH-1:0] in14,
  input [WIDTH-1:0] in15,
  input [WIDTH-1:0] in16,
  input [WIDTH-1:0] in17,
  input [WIDTH-1:0] in18,
  input [WIDTH-1:0] in19,
  input [WIDTH-1:0] in20,
  input [WIDTH-1:0] in21,
  input [WIDTH-1:0] in22,
  input [WIDTH-1:0] in23,
  input [WIDTH-1:0] in24,
  input [WIDTH-1:0] in25,
  input [WIDTH-1:0] in26,
  input [WIDTH-1:0] in27,
  input [WIDTH-1:0] in28,
  input [WIDTH-1:0] in29,
  input [WIDTH-1:0] in30,
  input [WIDTH-1:0] in31,
  input [WIDTH-1:0] in32,
  input [WIDTH-1:0] in33,
  input [WIDTH-1:0] in34,
  input [WIDTH-1:0] in35,
  input [WIDTH-1:0] in36,
  input [WIDTH-1:0] in37,
  input [WIDTH-1:0] in38,
  input [WIDTH-1:0] in39,
  input [WIDTH-1:0] in40,
  input [WIDTH-1:0] in41,
  input [WIDTH-1:0] in42,
  input [WIDTH-1:0] in43,
  input [WIDTH-1:0] in44,
  input [WIDTH-1:0] in45,
  input [WIDTH-1:0] in46,
  input [WIDTH-1:0] in47,
  input [WIDTH-1:0] in48,
  input [WIDTH-1:0] in49,
  input [WIDTH-1:0] in50,
  input [WIDTH-1:0] in51,
  input [WIDTH-1:0] in52,
  input [WIDTH-1:0] in53,
  input [WIDTH-1:0] in54,
  input [WIDTH-1:0] in55,
  input [WIDTH-1:0] in56,
  input [WIDTH-1:0] in57,
  input [WIDTH-1:0] in58,
  input [WIDTH-1:0] in59,
  input [WIDTH-1:0] in60,
  input [WIDTH-1:0] in61,
  input [WIDTH-1:0] in62,
  input [WIDTH-1:0] in63,
  input [WIDTH-1:0] in64,
  input [WIDTH-1:0] in65,
  input [WIDTH-1:0] in66,
  input [WIDTH-1:0] in67,
  input [WIDTH-1:0] in68,
  input [WIDTH-1:0] in69,
  input [WIDTH-1:0] in70,
  input [WIDTH-1:0] in71,
  input [WIDTH-1:0] in72,
  input [WIDTH-1:0] in73,
  input [WIDTH-1:0] in74,
  input [WIDTH-1:0] in75,
  input [WIDTH-1:0] in76,
  input [WIDTH-1:0] in77,
  input [WIDTH-1:0] in78,
  input [WIDTH-1:0] in79,
  input [WIDTH-1:0] in80,
  input [WIDTH-1:0] in81,
  input [WIDTH-1:0] in82,
  input [WIDTH-1:0] in83,
  input [WIDTH-1:0] in84,
  input [WIDTH-1:0] in85,
  input [WIDTH-1:0] in86,
  input [WIDTH-1:0] in87,
  input [WIDTH-1:0] in88,
  input [WIDTH-1:0] in89,
  input [WIDTH-1:0] in90,
  input [WIDTH-1:0] in91,
  input [WIDTH-1:0] in92,
  input [WIDTH-1:0] in93,
  input [WIDTH-1:0] in94,
  input [WIDTH-1:0] in95,
  input [WIDTH-1:0] in96,
  input [WIDTH-1:0] in97,
  input [WIDTH-1:0] in98,
  input [WIDTH-1:0] in99,
  input [WIDTH-1:0] in100,
  input [WIDTH-1:0] in101,
  input [WIDTH-1:0] in102,
  input [WIDTH-1:0] in103,
  input [WIDTH-1:0] in104,
  input [WIDTH-1:0] in105,
  input [WIDTH-1:0] in106,
  input [WIDTH-1:0] in107,
  input [WIDTH-1:0] in108,
  input [WIDTH-1:0] in109,
  input [WIDTH-1:0] in110,
  input [WIDTH-1:0] in111,
  input [WIDTH-1:0] in112,
  input [WIDTH-1:0] in113,
  input [WIDTH-1:0] in114,
  input [WIDTH-1:0] in115,
  input [WIDTH-1:0] in116,
  input [WIDTH-1:0] in117,
  input [WIDTH-1:0] in118,
  input [WIDTH-1:0] in119,
  input [WIDTH-1:0] in120,
  input [WIDTH-1:0] in121,
  input [WIDTH-1:0] in122,
  input [WIDTH-1:0] in123,
  input [WIDTH-1:0] in124,
  input [WIDTH-1:0] in125,
  input [WIDTH-1:0] in126,
  input [WIDTH-1:0] in127,
  output [WIDTH-1:0] out0,
  output [WIDTH-1:0] out1,
  output [WIDTH-1:0] out2,
  output [WIDTH-1:0] out3,
  output [WIDTH-1:0] out4,
  output [WIDTH-1:0] out5,
  output [WIDTH-1:0] out6,
  output [WIDTH-1:0] out7,
  output [WIDTH-1:0] out8,
  output [WIDTH-1:0] out9,
  output [WIDTH-1:0] out10,
  output [WIDTH-1:0] out11,
  output [WIDTH-1:0] out12,
  output [WIDTH-1:0] out13,
  output [WIDTH-1:0] out14,
  output [WIDTH-1:0] out15,
  output [WIDTH-1:0] out16,
  output [WIDTH-1:0] out17,
  output [WIDTH-1:0] out18,
  output [WIDTH-1:0] out19,
  output [WIDTH-1:0] out20,
  output [WIDTH-1:0] out21,
  output [WIDTH-1:0] out22,
  output [WIDTH-1:0] out23,
  output [WIDTH-1:0] out24,
  output [WIDTH-1:0] out25,
  output [WIDTH-1:0] out26,
  output [WIDTH-1:0] out27,
  output [WIDTH-1:0] out28,
  output [WIDTH-1:0] out29,
  output [WIDTH-1:0] out30,
  output [WIDTH-1:0] out31,
  output [WIDTH-1:0] out32,
  output [WIDTH-1:0] out33,
  output [WIDTH-1:0] out34,
  output [WIDTH-1:0] out35,
  output [WIDTH-1:0] out36,
  output [WIDTH-1:0] out37,
  output [WIDTH-1:0] out38,
  output [WIDTH-1:0] out39,
  output [WIDTH-1:0] out40,
  output [WIDTH-1:0] out41,
  output [WIDTH-1:0] out42,
  output [WIDTH-1:0] out43,
  output [WIDTH-1:0] out44,
  output [WIDTH-1:0] out45,
  output [WIDTH-1:0] out46,
  output [WIDTH-1:0] out47,
  output [WIDTH-1:0] out48,
  output [WIDTH-1:0] out49,
  output [WIDTH-1:0] out50,
  output [WIDTH-1:0] out51,
  output [WIDTH-1:0] out52,
  output [WIDTH-1:0] out53,
  output [WIDTH-1:0] out54,
  output [WIDTH-1:0] out55,
  output [WIDTH-1:0] out56,
  output [WIDTH-1:0] out57,
  output [WIDTH-1:0] out58,
  output [WIDTH-1:0] out59,
  output [WIDTH-1:0] out60,
  output [WIDTH-1:0] out61,
  output [WIDTH-1:0] out62,
  output [WIDTH-1:0] out63,
  output [WIDTH-1:0] out64,
  output [WIDTH-1:0] out65,
  output [WIDTH-1:0] out66,
  output [WIDTH-1:0] out67,
  output [WIDTH-1:0] out68,
  output [WIDTH-1:0] out69,
  output [WIDTH-1:0] out70,
  output [WIDTH-1:0] out71,
  output [WIDTH-1:0] out72,
  output [WIDTH-1:0] out73,
  output [WIDTH-1:0] out74,
  output [WIDTH-1:0] out75,
  output [WIDTH-1:0] out76,
  output [WIDTH-1:0] out77,
  output [WIDTH-1:0] out78,
  output [WIDTH-1:0] out79,
  output [WIDTH-1:0] out80,
  output [WIDTH-1:0] out81,
  output [WIDTH-1:0] out82,
  output [WIDTH-1:0] out83,
  output [WIDTH-1:0] out84,
  output [WIDTH-1:0] out85,
  output [WIDTH-1:0] out86,
  output [WIDTH-1:0] out87,
  output [WIDTH-1:0] out88,
  output [WIDTH-1:0] out89,
  output [WIDTH-1:0] out90,
  output [WIDTH-1:0] out91,
  output [WIDTH-1:0] out92,
  output [WIDTH-1:0] out93,
  output [WIDTH-1:0] out94,
  output [WIDTH-1:0] out95,
  output [WIDTH-1:0] out96,
  output [WIDTH-1:0] out97,
  output [WIDTH-1:0] out98,
  output [WIDTH-1:0] out99,
  output [WIDTH-1:0] out100,
  output [WIDTH-1:0] out101,
  output [WIDTH-1:0] out102,
  output [WIDTH-1:0] out103,
  output [WIDTH-1:0] out104,
  output [WIDTH-1:0] out105,
  output [WIDTH-1:0] out106,
  output [WIDTH-1:0] out107,
  output [WIDTH-1:0] out108,
  output [WIDTH-1:0] out109,
  output [WIDTH-1:0] out110,
  output [WIDTH-1:0] out111,
  output [WIDTH-1:0] out112,
  output [WIDTH-1:0] out113,
  output [WIDTH-1:0] out114,
  output [WIDTH-1:0] out115,
  output [WIDTH-1:0] out116,
  output [WIDTH-1:0] out117,
  output [WIDTH-1:0] out118,
  output [WIDTH-1:0] out119,
  output [WIDTH-1:0] out120,
  output [WIDTH-1:0] out121,
  output [WIDTH-1:0] out122,
  output [WIDTH-1:0] out123,
  output [WIDTH-1:0] out124,
  output [WIDTH-1:0] out125,
  output [WIDTH-1:0] out126,
  output [WIDTH-1:0] out127
);

  wire [1536-1:0] conf_out;
  wire [WIDTH-1:0] in_reg_wire_0 [0:128-1];
  wire [WIDTH-1:0] in_reg_wire_1 [0:128-1];
  wire [WIDTH-1:0] in_reg_wire_2 [0:128-1];
  wire [WIDTH-1:0] in_reg_wire_3 [0:128-1];
  wire [WIDTH-1:0] in_reg_wire_4 [0:128-1];
  wire [WIDTH-1:0] in_reg_wire_5 [0:128-1];
  wire [WIDTH-1:0] in_reg_wire_6 [0:128-1];
  wire [WIDTH-1:0] in_reg_wire_7 [0:128-1];
  wire [64-1:0] net_conf_bus [0:64-1];

  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg0
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus_in),
    .out(net_conf_bus[0])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(1),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_0
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[0]),
    .swicth_conf_out(conf_out[23:0])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg1
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[0]),
    .out(net_conf_bus[1])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(2),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_1
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[1]),
    .swicth_conf_out(conf_out[47:24])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg2
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[1]),
    .out(net_conf_bus[2])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(3),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_2
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[2]),
    .swicth_conf_out(conf_out[71:48])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg3
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[2]),
    .out(net_conf_bus[3])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(4),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_3
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[3]),
    .swicth_conf_out(conf_out[95:72])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg4
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[3]),
    .out(net_conf_bus[4])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(5),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_4
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[4]),
    .swicth_conf_out(conf_out[119:96])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg5
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[4]),
    .out(net_conf_bus[5])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(6),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_5
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[5]),
    .swicth_conf_out(conf_out[143:120])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg6
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[5]),
    .out(net_conf_bus[6])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(7),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_6
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[6]),
    .swicth_conf_out(conf_out[167:144])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg7
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[6]),
    .out(net_conf_bus[7])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(8),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_7
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[7]),
    .swicth_conf_out(conf_out[191:168])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg8
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[7]),
    .out(net_conf_bus[8])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(9),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_8
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[8]),
    .swicth_conf_out(conf_out[215:192])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg9
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[8]),
    .out(net_conf_bus[9])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(10),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_9
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[9]),
    .swicth_conf_out(conf_out[239:216])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg10
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[9]),
    .out(net_conf_bus[10])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(11),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_10
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[10]),
    .swicth_conf_out(conf_out[263:240])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg11
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[10]),
    .out(net_conf_bus[11])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(12),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_11
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[11]),
    .swicth_conf_out(conf_out[287:264])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg12
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[11]),
    .out(net_conf_bus[12])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(13),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_12
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[12]),
    .swicth_conf_out(conf_out[311:288])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg13
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[12]),
    .out(net_conf_bus[13])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(14),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_13
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[13]),
    .swicth_conf_out(conf_out[335:312])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg14
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[13]),
    .out(net_conf_bus[14])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(15),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_14
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[14]),
    .swicth_conf_out(conf_out[359:336])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg15
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[14]),
    .out(net_conf_bus[15])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(16),
    .STAGE(PIPE_EXTRA + 1)
  )
  swicth_conf_control_15
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[15]),
    .swicth_conf_out(conf_out[383:360])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg16
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[15]),
    .out(net_conf_bus[16])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(17),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_16
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[16]),
    .swicth_conf_out(conf_out[407:384])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg17
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[16]),
    .out(net_conf_bus[17])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(18),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_17
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[17]),
    .swicth_conf_out(conf_out[431:408])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg18
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[17]),
    .out(net_conf_bus[18])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(19),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_18
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[18]),
    .swicth_conf_out(conf_out[455:432])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg19
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[18]),
    .out(net_conf_bus[19])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(20),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_19
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[19]),
    .swicth_conf_out(conf_out[479:456])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg20
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[19]),
    .out(net_conf_bus[20])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(21),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_20
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[20]),
    .swicth_conf_out(conf_out[503:480])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg21
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[20]),
    .out(net_conf_bus[21])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(22),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_21
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[21]),
    .swicth_conf_out(conf_out[527:504])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg22
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[21]),
    .out(net_conf_bus[22])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(23),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_22
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[22]),
    .swicth_conf_out(conf_out[551:528])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg23
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[22]),
    .out(net_conf_bus[23])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(24),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_23
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[23]),
    .swicth_conf_out(conf_out[575:552])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg24
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[23]),
    .out(net_conf_bus[24])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(25),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_24
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[24]),
    .swicth_conf_out(conf_out[599:576])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg25
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[24]),
    .out(net_conf_bus[25])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(26),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_25
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[25]),
    .swicth_conf_out(conf_out[623:600])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg26
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[25]),
    .out(net_conf_bus[26])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(27),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_26
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[26]),
    .swicth_conf_out(conf_out[647:624])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg27
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[26]),
    .out(net_conf_bus[27])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(28),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_27
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[27]),
    .swicth_conf_out(conf_out[671:648])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg28
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[27]),
    .out(net_conf_bus[28])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(29),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_28
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[28]),
    .swicth_conf_out(conf_out[695:672])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg29
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[28]),
    .out(net_conf_bus[29])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(30),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_29
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[29]),
    .swicth_conf_out(conf_out[719:696])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg30
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[29]),
    .out(net_conf_bus[30])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(31),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_30
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[30]),
    .swicth_conf_out(conf_out[743:720])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg31
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[30]),
    .out(net_conf_bus[31])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(32),
    .STAGE(PIPE_EXTRA + 2)
  )
  swicth_conf_control_31
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[31]),
    .swicth_conf_out(conf_out[767:744])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg32
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[31]),
    .out(net_conf_bus[32])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(33),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_32
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[32]),
    .swicth_conf_out(conf_out[791:768])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg33
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[32]),
    .out(net_conf_bus[33])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(34),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_33
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[33]),
    .swicth_conf_out(conf_out[815:792])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg34
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[33]),
    .out(net_conf_bus[34])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(35),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_34
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[34]),
    .swicth_conf_out(conf_out[839:816])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg35
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[34]),
    .out(net_conf_bus[35])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(36),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_35
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[35]),
    .swicth_conf_out(conf_out[863:840])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg36
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[35]),
    .out(net_conf_bus[36])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(37),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_36
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[36]),
    .swicth_conf_out(conf_out[887:864])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg37
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[36]),
    .out(net_conf_bus[37])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(38),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_37
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[37]),
    .swicth_conf_out(conf_out[911:888])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg38
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[37]),
    .out(net_conf_bus[38])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(39),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_38
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[38]),
    .swicth_conf_out(conf_out[935:912])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg39
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[38]),
    .out(net_conf_bus[39])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(40),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_39
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[39]),
    .swicth_conf_out(conf_out[959:936])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg40
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[39]),
    .out(net_conf_bus[40])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(41),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_40
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[40]),
    .swicth_conf_out(conf_out[983:960])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg41
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[40]),
    .out(net_conf_bus[41])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(42),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_41
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[41]),
    .swicth_conf_out(conf_out[1007:984])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg42
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[41]),
    .out(net_conf_bus[42])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(43),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_42
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[42]),
    .swicth_conf_out(conf_out[1031:1008])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg43
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[42]),
    .out(net_conf_bus[43])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(44),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_43
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[43]),
    .swicth_conf_out(conf_out[1055:1032])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg44
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[43]),
    .out(net_conf_bus[44])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(45),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_44
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[44]),
    .swicth_conf_out(conf_out[1079:1056])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg45
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[44]),
    .out(net_conf_bus[45])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(46),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_45
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[45]),
    .swicth_conf_out(conf_out[1103:1080])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg46
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[45]),
    .out(net_conf_bus[46])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(47),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_46
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[46]),
    .swicth_conf_out(conf_out[1127:1104])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg47
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[46]),
    .out(net_conf_bus[47])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(48),
    .STAGE(PIPE_EXTRA + 3)
  )
  swicth_conf_control_47
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[47]),
    .swicth_conf_out(conf_out[1151:1128])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg48
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[47]),
    .out(net_conf_bus[48])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(49),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_48
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[48]),
    .swicth_conf_out(conf_out[1175:1152])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg49
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[48]),
    .out(net_conf_bus[49])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(50),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_49
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[49]),
    .swicth_conf_out(conf_out[1199:1176])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg50
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[49]),
    .out(net_conf_bus[50])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(51),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_50
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[50]),
    .swicth_conf_out(conf_out[1223:1200])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg51
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[50]),
    .out(net_conf_bus[51])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(52),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_51
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[51]),
    .swicth_conf_out(conf_out[1247:1224])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg52
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[51]),
    .out(net_conf_bus[52])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(53),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_52
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[52]),
    .swicth_conf_out(conf_out[1271:1248])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg53
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[52]),
    .out(net_conf_bus[53])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(54),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_53
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[53]),
    .swicth_conf_out(conf_out[1295:1272])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg54
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[53]),
    .out(net_conf_bus[54])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(55),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_54
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[54]),
    .swicth_conf_out(conf_out[1319:1296])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg55
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[54]),
    .out(net_conf_bus[55])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(56),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_55
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[55]),
    .swicth_conf_out(conf_out[1343:1320])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg56
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[55]),
    .out(net_conf_bus[56])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(57),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_56
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[56]),
    .swicth_conf_out(conf_out[1367:1344])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg57
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[56]),
    .out(net_conf_bus[57])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(58),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_57
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[57]),
    .swicth_conf_out(conf_out[1391:1368])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg58
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[57]),
    .out(net_conf_bus[58])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(59),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_58
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[58]),
    .swicth_conf_out(conf_out[1415:1392])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg59
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[58]),
    .out(net_conf_bus[59])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(60),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_59
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[59]),
    .swicth_conf_out(conf_out[1439:1416])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg60
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[59]),
    .out(net_conf_bus[60])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(61),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_60
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[60]),
    .swicth_conf_out(conf_out[1463:1440])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg61
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[60]),
    .out(net_conf_bus[61])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(62),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_61
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[61]),
    .swicth_conf_out(conf_out[1487:1464])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg62
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[61]),
    .out(net_conf_bus[62])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(63),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_62
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[62]),
    .swicth_conf_out(conf_out[1511:1488])
  );


  reg_pipe
  #(
    .NUM_STAGES(1),
    .DATA_WIDTH(64)
  )
  net_conf_bus_reg63
  (
    .clk(clk),
    .rst(1'b0),
    .en(1'b1),
    .in(net_conf_bus[62]),
    .out(net_conf_bus[63])
  );


  swicth_conf_control_branch_24_1
  #(
    .SWICTH_NUMBER(64),
    .STAGE(PIPE_EXTRA + 4)
  )
  swicth_conf_control_63
  (
    .clk(clk),
    .rst(rst),
    .en_pc_net(en),
    .conf_bus_in(net_conf_bus[63]),
    .swicth_conf_out(conf_out[1535:1512])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_0
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in0),
    .out(in_reg_wire_0[0])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_1
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in1),
    .out(in_reg_wire_0[1])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_2
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in2),
    .out(in_reg_wire_0[2])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_3
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in3),
    .out(in_reg_wire_0[3])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_4
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in4),
    .out(in_reg_wire_0[4])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_5
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in5),
    .out(in_reg_wire_0[5])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_6
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in6),
    .out(in_reg_wire_0[6])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_7
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in7),
    .out(in_reg_wire_0[7])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_8
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in8),
    .out(in_reg_wire_0[8])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_9
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in9),
    .out(in_reg_wire_0[9])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_10
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in10),
    .out(in_reg_wire_0[10])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_11
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in11),
    .out(in_reg_wire_0[11])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_12
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in12),
    .out(in_reg_wire_0[12])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_13
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in13),
    .out(in_reg_wire_0[13])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_14
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in14),
    .out(in_reg_wire_0[14])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_15
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in15),
    .out(in_reg_wire_0[15])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_16
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in16),
    .out(in_reg_wire_0[16])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_17
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in17),
    .out(in_reg_wire_0[17])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_18
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in18),
    .out(in_reg_wire_0[18])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_19
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in19),
    .out(in_reg_wire_0[19])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_20
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in20),
    .out(in_reg_wire_0[20])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_21
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in21),
    .out(in_reg_wire_0[21])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_22
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in22),
    .out(in_reg_wire_0[22])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_23
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in23),
    .out(in_reg_wire_0[23])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_24
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in24),
    .out(in_reg_wire_0[24])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_25
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in25),
    .out(in_reg_wire_0[25])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_26
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in26),
    .out(in_reg_wire_0[26])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_27
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in27),
    .out(in_reg_wire_0[27])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_28
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in28),
    .out(in_reg_wire_0[28])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_29
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in29),
    .out(in_reg_wire_0[29])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_30
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in30),
    .out(in_reg_wire_0[30])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_31
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in31),
    .out(in_reg_wire_0[31])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_32
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in32),
    .out(in_reg_wire_0[32])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_33
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in33),
    .out(in_reg_wire_0[33])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_34
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in34),
    .out(in_reg_wire_0[34])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_35
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in35),
    .out(in_reg_wire_0[35])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_36
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in36),
    .out(in_reg_wire_0[36])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_37
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in37),
    .out(in_reg_wire_0[37])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_38
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in38),
    .out(in_reg_wire_0[38])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_39
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in39),
    .out(in_reg_wire_0[39])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_40
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in40),
    .out(in_reg_wire_0[40])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_41
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in41),
    .out(in_reg_wire_0[41])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_42
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in42),
    .out(in_reg_wire_0[42])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_43
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in43),
    .out(in_reg_wire_0[43])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_44
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in44),
    .out(in_reg_wire_0[44])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_45
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in45),
    .out(in_reg_wire_0[45])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_46
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in46),
    .out(in_reg_wire_0[46])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_47
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in47),
    .out(in_reg_wire_0[47])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_48
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in48),
    .out(in_reg_wire_0[48])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_49
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in49),
    .out(in_reg_wire_0[49])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_50
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in50),
    .out(in_reg_wire_0[50])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_51
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in51),
    .out(in_reg_wire_0[51])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_52
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in52),
    .out(in_reg_wire_0[52])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_53
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in53),
    .out(in_reg_wire_0[53])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_54
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in54),
    .out(in_reg_wire_0[54])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_55
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in55),
    .out(in_reg_wire_0[55])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_56
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in56),
    .out(in_reg_wire_0[56])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_57
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in57),
    .out(in_reg_wire_0[57])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_58
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in58),
    .out(in_reg_wire_0[58])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_59
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in59),
    .out(in_reg_wire_0[59])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_60
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in60),
    .out(in_reg_wire_0[60])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_61
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in61),
    .out(in_reg_wire_0[61])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_62
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in62),
    .out(in_reg_wire_0[62])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_63
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in63),
    .out(in_reg_wire_0[63])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_64
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in64),
    .out(in_reg_wire_0[64])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_65
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in65),
    .out(in_reg_wire_0[65])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_66
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in66),
    .out(in_reg_wire_0[66])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_67
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in67),
    .out(in_reg_wire_0[67])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_68
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in68),
    .out(in_reg_wire_0[68])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_69
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in69),
    .out(in_reg_wire_0[69])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_70
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in70),
    .out(in_reg_wire_0[70])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_71
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in71),
    .out(in_reg_wire_0[71])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_72
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in72),
    .out(in_reg_wire_0[72])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_73
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in73),
    .out(in_reg_wire_0[73])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_74
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in74),
    .out(in_reg_wire_0[74])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_75
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in75),
    .out(in_reg_wire_0[75])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_76
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in76),
    .out(in_reg_wire_0[76])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_77
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in77),
    .out(in_reg_wire_0[77])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_78
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in78),
    .out(in_reg_wire_0[78])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_79
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in79),
    .out(in_reg_wire_0[79])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_80
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in80),
    .out(in_reg_wire_0[80])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_81
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in81),
    .out(in_reg_wire_0[81])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_82
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in82),
    .out(in_reg_wire_0[82])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_83
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in83),
    .out(in_reg_wire_0[83])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_84
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in84),
    .out(in_reg_wire_0[84])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_85
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in85),
    .out(in_reg_wire_0[85])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_86
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in86),
    .out(in_reg_wire_0[86])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_87
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in87),
    .out(in_reg_wire_0[87])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_88
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in88),
    .out(in_reg_wire_0[88])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_89
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in89),
    .out(in_reg_wire_0[89])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_90
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in90),
    .out(in_reg_wire_0[90])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_91
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in91),
    .out(in_reg_wire_0[91])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_92
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in92),
    .out(in_reg_wire_0[92])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_93
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in93),
    .out(in_reg_wire_0[93])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_94
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in94),
    .out(in_reg_wire_0[94])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_95
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in95),
    .out(in_reg_wire_0[95])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_96
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in96),
    .out(in_reg_wire_0[96])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_97
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in97),
    .out(in_reg_wire_0[97])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_98
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in98),
    .out(in_reg_wire_0[98])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_99
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in99),
    .out(in_reg_wire_0[99])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_100
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in100),
    .out(in_reg_wire_0[100])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_101
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in101),
    .out(in_reg_wire_0[101])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_102
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in102),
    .out(in_reg_wire_0[102])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_103
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in103),
    .out(in_reg_wire_0[103])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_104
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in104),
    .out(in_reg_wire_0[104])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_105
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in105),
    .out(in_reg_wire_0[105])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_106
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in106),
    .out(in_reg_wire_0[106])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_107
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in107),
    .out(in_reg_wire_0[107])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_108
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in108),
    .out(in_reg_wire_0[108])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_109
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in109),
    .out(in_reg_wire_0[109])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_110
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in110),
    .out(in_reg_wire_0[110])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_111
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in111),
    .out(in_reg_wire_0[111])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_112
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in112),
    .out(in_reg_wire_0[112])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_113
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in113),
    .out(in_reg_wire_0[113])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_114
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in114),
    .out(in_reg_wire_0[114])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_115
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in115),
    .out(in_reg_wire_0[115])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_116
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in116),
    .out(in_reg_wire_0[116])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_117
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in117),
    .out(in_reg_wire_0[117])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_118
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in118),
    .out(in_reg_wire_0[118])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_119
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in119),
    .out(in_reg_wire_0[119])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_120
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in120),
    .out(in_reg_wire_0[120])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_121
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in121),
    .out(in_reg_wire_0[121])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_122
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in122),
    .out(in_reg_wire_0[122])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_123
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in123),
    .out(in_reg_wire_0[123])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_124
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in124),
    .out(in_reg_wire_0[124])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_125
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in125),
    .out(in_reg_wire_0[125])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_126
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in126),
    .out(in_reg_wire_0[126])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_0_127
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in127),
    .out(in_reg_wire_0[127])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_0
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[0]),
    .out(in_reg_wire_2[0])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_1
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[1]),
    .out(in_reg_wire_2[1])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_2
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[2]),
    .out(in_reg_wire_2[2])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_3
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[3]),
    .out(in_reg_wire_2[3])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_4
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[4]),
    .out(in_reg_wire_2[4])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_5
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[5]),
    .out(in_reg_wire_2[5])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_6
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[6]),
    .out(in_reg_wire_2[6])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_7
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[7]),
    .out(in_reg_wire_2[7])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_8
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[8]),
    .out(in_reg_wire_2[8])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_9
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[9]),
    .out(in_reg_wire_2[9])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_10
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[10]),
    .out(in_reg_wire_2[10])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_11
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[11]),
    .out(in_reg_wire_2[11])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_12
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[12]),
    .out(in_reg_wire_2[12])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_13
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[13]),
    .out(in_reg_wire_2[13])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_14
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[14]),
    .out(in_reg_wire_2[14])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_15
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[15]),
    .out(in_reg_wire_2[15])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_16
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[16]),
    .out(in_reg_wire_2[16])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_17
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[17]),
    .out(in_reg_wire_2[17])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_18
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[18]),
    .out(in_reg_wire_2[18])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_19
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[19]),
    .out(in_reg_wire_2[19])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_20
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[20]),
    .out(in_reg_wire_2[20])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_21
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[21]),
    .out(in_reg_wire_2[21])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_22
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[22]),
    .out(in_reg_wire_2[22])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_23
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[23]),
    .out(in_reg_wire_2[23])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_24
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[24]),
    .out(in_reg_wire_2[24])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_25
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[25]),
    .out(in_reg_wire_2[25])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_26
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[26]),
    .out(in_reg_wire_2[26])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_27
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[27]),
    .out(in_reg_wire_2[27])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_28
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[28]),
    .out(in_reg_wire_2[28])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_29
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[29]),
    .out(in_reg_wire_2[29])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_30
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[30]),
    .out(in_reg_wire_2[30])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_31
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[31]),
    .out(in_reg_wire_2[31])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_32
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[32]),
    .out(in_reg_wire_2[32])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_33
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[33]),
    .out(in_reg_wire_2[33])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_34
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[34]),
    .out(in_reg_wire_2[34])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_35
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[35]),
    .out(in_reg_wire_2[35])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_36
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[36]),
    .out(in_reg_wire_2[36])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_37
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[37]),
    .out(in_reg_wire_2[37])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_38
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[38]),
    .out(in_reg_wire_2[38])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_39
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[39]),
    .out(in_reg_wire_2[39])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_40
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[40]),
    .out(in_reg_wire_2[40])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_41
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[41]),
    .out(in_reg_wire_2[41])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_42
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[42]),
    .out(in_reg_wire_2[42])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_43
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[43]),
    .out(in_reg_wire_2[43])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_44
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[44]),
    .out(in_reg_wire_2[44])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_45
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[45]),
    .out(in_reg_wire_2[45])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_46
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[46]),
    .out(in_reg_wire_2[46])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_47
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[47]),
    .out(in_reg_wire_2[47])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_48
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[48]),
    .out(in_reg_wire_2[48])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_49
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[49]),
    .out(in_reg_wire_2[49])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_50
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[50]),
    .out(in_reg_wire_2[50])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_51
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[51]),
    .out(in_reg_wire_2[51])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_52
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[52]),
    .out(in_reg_wire_2[52])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_53
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[53]),
    .out(in_reg_wire_2[53])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_54
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[54]),
    .out(in_reg_wire_2[54])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_55
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[55]),
    .out(in_reg_wire_2[55])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_56
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[56]),
    .out(in_reg_wire_2[56])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_57
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[57]),
    .out(in_reg_wire_2[57])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_58
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[58]),
    .out(in_reg_wire_2[58])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_59
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[59]),
    .out(in_reg_wire_2[59])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_60
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[60]),
    .out(in_reg_wire_2[60])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_61
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[61]),
    .out(in_reg_wire_2[61])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_62
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[62]),
    .out(in_reg_wire_2[62])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_63
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[63]),
    .out(in_reg_wire_2[63])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_64
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[64]),
    .out(in_reg_wire_2[64])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_65
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[65]),
    .out(in_reg_wire_2[65])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_66
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[66]),
    .out(in_reg_wire_2[66])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_67
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[67]),
    .out(in_reg_wire_2[67])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_68
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[68]),
    .out(in_reg_wire_2[68])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_69
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[69]),
    .out(in_reg_wire_2[69])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_70
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[70]),
    .out(in_reg_wire_2[70])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_71
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[71]),
    .out(in_reg_wire_2[71])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_72
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[72]),
    .out(in_reg_wire_2[72])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_73
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[73]),
    .out(in_reg_wire_2[73])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_74
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[74]),
    .out(in_reg_wire_2[74])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_75
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[75]),
    .out(in_reg_wire_2[75])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_76
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[76]),
    .out(in_reg_wire_2[76])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_77
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[77]),
    .out(in_reg_wire_2[77])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_78
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[78]),
    .out(in_reg_wire_2[78])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_79
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[79]),
    .out(in_reg_wire_2[79])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_80
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[80]),
    .out(in_reg_wire_2[80])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_81
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[81]),
    .out(in_reg_wire_2[81])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_82
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[82]),
    .out(in_reg_wire_2[82])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_83
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[83]),
    .out(in_reg_wire_2[83])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_84
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[84]),
    .out(in_reg_wire_2[84])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_85
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[85]),
    .out(in_reg_wire_2[85])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_86
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[86]),
    .out(in_reg_wire_2[86])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_87
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[87]),
    .out(in_reg_wire_2[87])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_88
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[88]),
    .out(in_reg_wire_2[88])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_89
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[89]),
    .out(in_reg_wire_2[89])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_90
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[90]),
    .out(in_reg_wire_2[90])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_91
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[91]),
    .out(in_reg_wire_2[91])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_92
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[92]),
    .out(in_reg_wire_2[92])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_93
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[93]),
    .out(in_reg_wire_2[93])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_94
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[94]),
    .out(in_reg_wire_2[94])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_95
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[95]),
    .out(in_reg_wire_2[95])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_96
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[96]),
    .out(in_reg_wire_2[96])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_97
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[97]),
    .out(in_reg_wire_2[97])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_98
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[98]),
    .out(in_reg_wire_2[98])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_99
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[99]),
    .out(in_reg_wire_2[99])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_100
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[100]),
    .out(in_reg_wire_2[100])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_101
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[101]),
    .out(in_reg_wire_2[101])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_102
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[102]),
    .out(in_reg_wire_2[102])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_103
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[103]),
    .out(in_reg_wire_2[103])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_104
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[104]),
    .out(in_reg_wire_2[104])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_105
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[105]),
    .out(in_reg_wire_2[105])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_106
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[106]),
    .out(in_reg_wire_2[106])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_107
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[107]),
    .out(in_reg_wire_2[107])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_108
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[108]),
    .out(in_reg_wire_2[108])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_109
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[109]),
    .out(in_reg_wire_2[109])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_110
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[110]),
    .out(in_reg_wire_2[110])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_111
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[111]),
    .out(in_reg_wire_2[111])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_112
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[112]),
    .out(in_reg_wire_2[112])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_113
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[113]),
    .out(in_reg_wire_2[113])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_114
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[114]),
    .out(in_reg_wire_2[114])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_115
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[115]),
    .out(in_reg_wire_2[115])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_116
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[116]),
    .out(in_reg_wire_2[116])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_117
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[117]),
    .out(in_reg_wire_2[117])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_118
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[118]),
    .out(in_reg_wire_2[118])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_119
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[119]),
    .out(in_reg_wire_2[119])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_120
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[120]),
    .out(in_reg_wire_2[120])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_121
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[121]),
    .out(in_reg_wire_2[121])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_122
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[122]),
    .out(in_reg_wire_2[122])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_123
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[123]),
    .out(in_reg_wire_2[123])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_124
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[124]),
    .out(in_reg_wire_2[124])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_125
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[125]),
    .out(in_reg_wire_2[125])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_126
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[126]),
    .out(in_reg_wire_2[126])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_1_127
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_1[127]),
    .out(in_reg_wire_2[127])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_0
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[0]),
    .out(in_reg_wire_4[0])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_1
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[1]),
    .out(in_reg_wire_4[1])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_2
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[2]),
    .out(in_reg_wire_4[2])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_3
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[3]),
    .out(in_reg_wire_4[3])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_4
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[4]),
    .out(in_reg_wire_4[4])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_5
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[5]),
    .out(in_reg_wire_4[5])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_6
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[6]),
    .out(in_reg_wire_4[6])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_7
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[7]),
    .out(in_reg_wire_4[7])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_8
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[8]),
    .out(in_reg_wire_4[8])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_9
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[9]),
    .out(in_reg_wire_4[9])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_10
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[10]),
    .out(in_reg_wire_4[10])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_11
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[11]),
    .out(in_reg_wire_4[11])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_12
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[12]),
    .out(in_reg_wire_4[12])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_13
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[13]),
    .out(in_reg_wire_4[13])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_14
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[14]),
    .out(in_reg_wire_4[14])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_15
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[15]),
    .out(in_reg_wire_4[15])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_16
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[16]),
    .out(in_reg_wire_4[16])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_17
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[17]),
    .out(in_reg_wire_4[17])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_18
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[18]),
    .out(in_reg_wire_4[18])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_19
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[19]),
    .out(in_reg_wire_4[19])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_20
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[20]),
    .out(in_reg_wire_4[20])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_21
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[21]),
    .out(in_reg_wire_4[21])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_22
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[22]),
    .out(in_reg_wire_4[22])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_23
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[23]),
    .out(in_reg_wire_4[23])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_24
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[24]),
    .out(in_reg_wire_4[24])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_25
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[25]),
    .out(in_reg_wire_4[25])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_26
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[26]),
    .out(in_reg_wire_4[26])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_27
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[27]),
    .out(in_reg_wire_4[27])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_28
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[28]),
    .out(in_reg_wire_4[28])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_29
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[29]),
    .out(in_reg_wire_4[29])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_30
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[30]),
    .out(in_reg_wire_4[30])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_31
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[31]),
    .out(in_reg_wire_4[31])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_32
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[32]),
    .out(in_reg_wire_4[32])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_33
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[33]),
    .out(in_reg_wire_4[33])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_34
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[34]),
    .out(in_reg_wire_4[34])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_35
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[35]),
    .out(in_reg_wire_4[35])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_36
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[36]),
    .out(in_reg_wire_4[36])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_37
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[37]),
    .out(in_reg_wire_4[37])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_38
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[38]),
    .out(in_reg_wire_4[38])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_39
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[39]),
    .out(in_reg_wire_4[39])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_40
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[40]),
    .out(in_reg_wire_4[40])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_41
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[41]),
    .out(in_reg_wire_4[41])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_42
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[42]),
    .out(in_reg_wire_4[42])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_43
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[43]),
    .out(in_reg_wire_4[43])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_44
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[44]),
    .out(in_reg_wire_4[44])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_45
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[45]),
    .out(in_reg_wire_4[45])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_46
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[46]),
    .out(in_reg_wire_4[46])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_47
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[47]),
    .out(in_reg_wire_4[47])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_48
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[48]),
    .out(in_reg_wire_4[48])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_49
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[49]),
    .out(in_reg_wire_4[49])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_50
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[50]),
    .out(in_reg_wire_4[50])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_51
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[51]),
    .out(in_reg_wire_4[51])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_52
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[52]),
    .out(in_reg_wire_4[52])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_53
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[53]),
    .out(in_reg_wire_4[53])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_54
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[54]),
    .out(in_reg_wire_4[54])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_55
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[55]),
    .out(in_reg_wire_4[55])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_56
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[56]),
    .out(in_reg_wire_4[56])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_57
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[57]),
    .out(in_reg_wire_4[57])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_58
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[58]),
    .out(in_reg_wire_4[58])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_59
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[59]),
    .out(in_reg_wire_4[59])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_60
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[60]),
    .out(in_reg_wire_4[60])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_61
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[61]),
    .out(in_reg_wire_4[61])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_62
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[62]),
    .out(in_reg_wire_4[62])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_63
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[63]),
    .out(in_reg_wire_4[63])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_64
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[64]),
    .out(in_reg_wire_4[64])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_65
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[65]),
    .out(in_reg_wire_4[65])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_66
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[66]),
    .out(in_reg_wire_4[66])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_67
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[67]),
    .out(in_reg_wire_4[67])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_68
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[68]),
    .out(in_reg_wire_4[68])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_69
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[69]),
    .out(in_reg_wire_4[69])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_70
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[70]),
    .out(in_reg_wire_4[70])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_71
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[71]),
    .out(in_reg_wire_4[71])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_72
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[72]),
    .out(in_reg_wire_4[72])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_73
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[73]),
    .out(in_reg_wire_4[73])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_74
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[74]),
    .out(in_reg_wire_4[74])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_75
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[75]),
    .out(in_reg_wire_4[75])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_76
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[76]),
    .out(in_reg_wire_4[76])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_77
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[77]),
    .out(in_reg_wire_4[77])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_78
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[78]),
    .out(in_reg_wire_4[78])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_79
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[79]),
    .out(in_reg_wire_4[79])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_80
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[80]),
    .out(in_reg_wire_4[80])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_81
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[81]),
    .out(in_reg_wire_4[81])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_82
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[82]),
    .out(in_reg_wire_4[82])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_83
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[83]),
    .out(in_reg_wire_4[83])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_84
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[84]),
    .out(in_reg_wire_4[84])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_85
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[85]),
    .out(in_reg_wire_4[85])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_86
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[86]),
    .out(in_reg_wire_4[86])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_87
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[87]),
    .out(in_reg_wire_4[87])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_88
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[88]),
    .out(in_reg_wire_4[88])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_89
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[89]),
    .out(in_reg_wire_4[89])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_90
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[90]),
    .out(in_reg_wire_4[90])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_91
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[91]),
    .out(in_reg_wire_4[91])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_92
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[92]),
    .out(in_reg_wire_4[92])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_93
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[93]),
    .out(in_reg_wire_4[93])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_94
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[94]),
    .out(in_reg_wire_4[94])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_95
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[95]),
    .out(in_reg_wire_4[95])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_96
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[96]),
    .out(in_reg_wire_4[96])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_97
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[97]),
    .out(in_reg_wire_4[97])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_98
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[98]),
    .out(in_reg_wire_4[98])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_99
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[99]),
    .out(in_reg_wire_4[99])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_100
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[100]),
    .out(in_reg_wire_4[100])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_101
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[101]),
    .out(in_reg_wire_4[101])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_102
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[102]),
    .out(in_reg_wire_4[102])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_103
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[103]),
    .out(in_reg_wire_4[103])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_104
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[104]),
    .out(in_reg_wire_4[104])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_105
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[105]),
    .out(in_reg_wire_4[105])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_106
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[106]),
    .out(in_reg_wire_4[106])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_107
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[107]),
    .out(in_reg_wire_4[107])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_108
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[108]),
    .out(in_reg_wire_4[108])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_109
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[109]),
    .out(in_reg_wire_4[109])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_110
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[110]),
    .out(in_reg_wire_4[110])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_111
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[111]),
    .out(in_reg_wire_4[111])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_112
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[112]),
    .out(in_reg_wire_4[112])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_113
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[113]),
    .out(in_reg_wire_4[113])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_114
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[114]),
    .out(in_reg_wire_4[114])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_115
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[115]),
    .out(in_reg_wire_4[115])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_116
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[116]),
    .out(in_reg_wire_4[116])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_117
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[117]),
    .out(in_reg_wire_4[117])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_118
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[118]),
    .out(in_reg_wire_4[118])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_119
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[119]),
    .out(in_reg_wire_4[119])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_120
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[120]),
    .out(in_reg_wire_4[120])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_121
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[121]),
    .out(in_reg_wire_4[121])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_122
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[122]),
    .out(in_reg_wire_4[122])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_123
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[123]),
    .out(in_reg_wire_4[123])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_124
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[124]),
    .out(in_reg_wire_4[124])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_125
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[125]),
    .out(in_reg_wire_4[125])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_126
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[126]),
    .out(in_reg_wire_4[126])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_2_127
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_3[127]),
    .out(in_reg_wire_4[127])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_0
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[0]),
    .out(in_reg_wire_6[0])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_1
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[1]),
    .out(in_reg_wire_6[1])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_2
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[2]),
    .out(in_reg_wire_6[2])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_3
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[3]),
    .out(in_reg_wire_6[3])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_4
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[4]),
    .out(in_reg_wire_6[4])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_5
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[5]),
    .out(in_reg_wire_6[5])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_6
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[6]),
    .out(in_reg_wire_6[6])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_7
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[7]),
    .out(in_reg_wire_6[7])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_8
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[8]),
    .out(in_reg_wire_6[8])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_9
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[9]),
    .out(in_reg_wire_6[9])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_10
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[10]),
    .out(in_reg_wire_6[10])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_11
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[11]),
    .out(in_reg_wire_6[11])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_12
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[12]),
    .out(in_reg_wire_6[12])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_13
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[13]),
    .out(in_reg_wire_6[13])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_14
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[14]),
    .out(in_reg_wire_6[14])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_15
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[15]),
    .out(in_reg_wire_6[15])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_16
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[16]),
    .out(in_reg_wire_6[16])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_17
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[17]),
    .out(in_reg_wire_6[17])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_18
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[18]),
    .out(in_reg_wire_6[18])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_19
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[19]),
    .out(in_reg_wire_6[19])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_20
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[20]),
    .out(in_reg_wire_6[20])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_21
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[21]),
    .out(in_reg_wire_6[21])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_22
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[22]),
    .out(in_reg_wire_6[22])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_23
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[23]),
    .out(in_reg_wire_6[23])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_24
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[24]),
    .out(in_reg_wire_6[24])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_25
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[25]),
    .out(in_reg_wire_6[25])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_26
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[26]),
    .out(in_reg_wire_6[26])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_27
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[27]),
    .out(in_reg_wire_6[27])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_28
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[28]),
    .out(in_reg_wire_6[28])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_29
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[29]),
    .out(in_reg_wire_6[29])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_30
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[30]),
    .out(in_reg_wire_6[30])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_31
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[31]),
    .out(in_reg_wire_6[31])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_32
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[32]),
    .out(in_reg_wire_6[32])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_33
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[33]),
    .out(in_reg_wire_6[33])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_34
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[34]),
    .out(in_reg_wire_6[34])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_35
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[35]),
    .out(in_reg_wire_6[35])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_36
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[36]),
    .out(in_reg_wire_6[36])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_37
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[37]),
    .out(in_reg_wire_6[37])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_38
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[38]),
    .out(in_reg_wire_6[38])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_39
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[39]),
    .out(in_reg_wire_6[39])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_40
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[40]),
    .out(in_reg_wire_6[40])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_41
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[41]),
    .out(in_reg_wire_6[41])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_42
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[42]),
    .out(in_reg_wire_6[42])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_43
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[43]),
    .out(in_reg_wire_6[43])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_44
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[44]),
    .out(in_reg_wire_6[44])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_45
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[45]),
    .out(in_reg_wire_6[45])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_46
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[46]),
    .out(in_reg_wire_6[46])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_47
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[47]),
    .out(in_reg_wire_6[47])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_48
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[48]),
    .out(in_reg_wire_6[48])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_49
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[49]),
    .out(in_reg_wire_6[49])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_50
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[50]),
    .out(in_reg_wire_6[50])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_51
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[51]),
    .out(in_reg_wire_6[51])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_52
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[52]),
    .out(in_reg_wire_6[52])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_53
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[53]),
    .out(in_reg_wire_6[53])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_54
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[54]),
    .out(in_reg_wire_6[54])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_55
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[55]),
    .out(in_reg_wire_6[55])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_56
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[56]),
    .out(in_reg_wire_6[56])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_57
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[57]),
    .out(in_reg_wire_6[57])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_58
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[58]),
    .out(in_reg_wire_6[58])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_59
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[59]),
    .out(in_reg_wire_6[59])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_60
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[60]),
    .out(in_reg_wire_6[60])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_61
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[61]),
    .out(in_reg_wire_6[61])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_62
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[62]),
    .out(in_reg_wire_6[62])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_63
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[63]),
    .out(in_reg_wire_6[63])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_64
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[64]),
    .out(in_reg_wire_6[64])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_65
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[65]),
    .out(in_reg_wire_6[65])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_66
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[66]),
    .out(in_reg_wire_6[66])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_67
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[67]),
    .out(in_reg_wire_6[67])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_68
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[68]),
    .out(in_reg_wire_6[68])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_69
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[69]),
    .out(in_reg_wire_6[69])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_70
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[70]),
    .out(in_reg_wire_6[70])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_71
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[71]),
    .out(in_reg_wire_6[71])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_72
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[72]),
    .out(in_reg_wire_6[72])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_73
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[73]),
    .out(in_reg_wire_6[73])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_74
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[74]),
    .out(in_reg_wire_6[74])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_75
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[75]),
    .out(in_reg_wire_6[75])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_76
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[76]),
    .out(in_reg_wire_6[76])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_77
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[77]),
    .out(in_reg_wire_6[77])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_78
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[78]),
    .out(in_reg_wire_6[78])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_79
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[79]),
    .out(in_reg_wire_6[79])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_80
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[80]),
    .out(in_reg_wire_6[80])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_81
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[81]),
    .out(in_reg_wire_6[81])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_82
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[82]),
    .out(in_reg_wire_6[82])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_83
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[83]),
    .out(in_reg_wire_6[83])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_84
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[84]),
    .out(in_reg_wire_6[84])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_85
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[85]),
    .out(in_reg_wire_6[85])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_86
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[86]),
    .out(in_reg_wire_6[86])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_87
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[87]),
    .out(in_reg_wire_6[87])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_88
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[88]),
    .out(in_reg_wire_6[88])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_89
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[89]),
    .out(in_reg_wire_6[89])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_90
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[90]),
    .out(in_reg_wire_6[90])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_91
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[91]),
    .out(in_reg_wire_6[91])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_92
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[92]),
    .out(in_reg_wire_6[92])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_93
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[93]),
    .out(in_reg_wire_6[93])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_94
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[94]),
    .out(in_reg_wire_6[94])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_95
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[95]),
    .out(in_reg_wire_6[95])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_96
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[96]),
    .out(in_reg_wire_6[96])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_97
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[97]),
    .out(in_reg_wire_6[97])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_98
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[98]),
    .out(in_reg_wire_6[98])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_99
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[99]),
    .out(in_reg_wire_6[99])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_100
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[100]),
    .out(in_reg_wire_6[100])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_101
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[101]),
    .out(in_reg_wire_6[101])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_102
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[102]),
    .out(in_reg_wire_6[102])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_103
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[103]),
    .out(in_reg_wire_6[103])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_104
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[104]),
    .out(in_reg_wire_6[104])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_105
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[105]),
    .out(in_reg_wire_6[105])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_106
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[106]),
    .out(in_reg_wire_6[106])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_107
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[107]),
    .out(in_reg_wire_6[107])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_108
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[108]),
    .out(in_reg_wire_6[108])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_109
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[109]),
    .out(in_reg_wire_6[109])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_110
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[110]),
    .out(in_reg_wire_6[110])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_111
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[111]),
    .out(in_reg_wire_6[111])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_112
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[112]),
    .out(in_reg_wire_6[112])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_113
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[113]),
    .out(in_reg_wire_6[113])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_114
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[114]),
    .out(in_reg_wire_6[114])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_115
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[115]),
    .out(in_reg_wire_6[115])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_116
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[116]),
    .out(in_reg_wire_6[116])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_117
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[117]),
    .out(in_reg_wire_6[117])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_118
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[118]),
    .out(in_reg_wire_6[118])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_119
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[119]),
    .out(in_reg_wire_6[119])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_120
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[120]),
    .out(in_reg_wire_6[120])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_121
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[121]),
    .out(in_reg_wire_6[121])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_122
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[122]),
    .out(in_reg_wire_6[122])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_123
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[123]),
    .out(in_reg_wire_6[123])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_124
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[124]),
    .out(in_reg_wire_6[124])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_125
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[125]),
    .out(in_reg_wire_6[125])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_126
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[126]),
    .out(in_reg_wire_6[126])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_3_127
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_5[127]),
    .out(in_reg_wire_6[127])
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_0
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[0]),
    .out(out0)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_1
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[1]),
    .out(out8)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_2
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[2]),
    .out(out16)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_3
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[3]),
    .out(out24)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_4
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[4]),
    .out(out32)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_5
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[5]),
    .out(out40)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_6
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[6]),
    .out(out48)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_7
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[7]),
    .out(out56)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_8
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[8]),
    .out(out64)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_9
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[9]),
    .out(out72)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_10
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[10]),
    .out(out80)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_11
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[11]),
    .out(out88)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_12
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[12]),
    .out(out96)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_13
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[13]),
    .out(out104)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_14
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[14]),
    .out(out112)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_15
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[15]),
    .out(out120)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_16
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[16]),
    .out(out1)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_17
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[17]),
    .out(out9)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_18
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[18]),
    .out(out17)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_19
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[19]),
    .out(out25)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_20
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[20]),
    .out(out33)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_21
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[21]),
    .out(out41)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_22
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[22]),
    .out(out49)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_23
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[23]),
    .out(out57)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_24
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[24]),
    .out(out65)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_25
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[25]),
    .out(out73)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_26
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[26]),
    .out(out81)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_27
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[27]),
    .out(out89)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_28
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[28]),
    .out(out97)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_29
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[29]),
    .out(out105)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_30
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[30]),
    .out(out113)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_31
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[31]),
    .out(out121)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_32
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[32]),
    .out(out2)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_33
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[33]),
    .out(out10)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_34
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[34]),
    .out(out18)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_35
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[35]),
    .out(out26)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_36
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[36]),
    .out(out34)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_37
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[37]),
    .out(out42)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_38
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[38]),
    .out(out50)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_39
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[39]),
    .out(out58)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_40
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[40]),
    .out(out66)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_41
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[41]),
    .out(out74)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_42
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[42]),
    .out(out82)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_43
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[43]),
    .out(out90)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_44
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[44]),
    .out(out98)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_45
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[45]),
    .out(out106)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_46
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[46]),
    .out(out114)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_47
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[47]),
    .out(out122)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_48
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[48]),
    .out(out3)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_49
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[49]),
    .out(out11)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_50
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[50]),
    .out(out19)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_51
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[51]),
    .out(out27)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_52
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[52]),
    .out(out35)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_53
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[53]),
    .out(out43)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_54
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[54]),
    .out(out51)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_55
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[55]),
    .out(out59)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_56
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[56]),
    .out(out67)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_57
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[57]),
    .out(out75)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_58
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[58]),
    .out(out83)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_59
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[59]),
    .out(out91)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_60
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[60]),
    .out(out99)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_61
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[61]),
    .out(out107)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_62
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[62]),
    .out(out115)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_63
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[63]),
    .out(out123)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_64
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[64]),
    .out(out4)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_65
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[65]),
    .out(out12)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_66
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[66]),
    .out(out20)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_67
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[67]),
    .out(out28)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_68
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[68]),
    .out(out36)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_69
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[69]),
    .out(out44)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_70
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[70]),
    .out(out52)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_71
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[71]),
    .out(out60)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_72
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[72]),
    .out(out68)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_73
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[73]),
    .out(out76)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_74
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[74]),
    .out(out84)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_75
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[75]),
    .out(out92)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_76
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[76]),
    .out(out100)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_77
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[77]),
    .out(out108)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_78
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[78]),
    .out(out116)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_79
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[79]),
    .out(out124)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_80
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[80]),
    .out(out5)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_81
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[81]),
    .out(out13)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_82
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[82]),
    .out(out21)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_83
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[83]),
    .out(out29)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_84
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[84]),
    .out(out37)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_85
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[85]),
    .out(out45)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_86
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[86]),
    .out(out53)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_87
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[87]),
    .out(out61)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_88
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[88]),
    .out(out69)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_89
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[89]),
    .out(out77)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_90
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[90]),
    .out(out85)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_91
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[91]),
    .out(out93)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_92
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[92]),
    .out(out101)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_93
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[93]),
    .out(out109)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_94
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[94]),
    .out(out117)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_95
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[95]),
    .out(out125)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_96
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[96]),
    .out(out6)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_97
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[97]),
    .out(out14)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_98
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[98]),
    .out(out22)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_99
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[99]),
    .out(out30)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_100
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[100]),
    .out(out38)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_101
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[101]),
    .out(out46)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_102
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[102]),
    .out(out54)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_103
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[103]),
    .out(out62)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_104
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[104]),
    .out(out70)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_105
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[105]),
    .out(out78)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_106
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[106]),
    .out(out86)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_107
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[107]),
    .out(out94)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_108
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[108]),
    .out(out102)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_109
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[109]),
    .out(out110)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_110
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[110]),
    .out(out118)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_111
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[111]),
    .out(out126)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_112
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[112]),
    .out(out7)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_113
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[113]),
    .out(out15)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_114
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[114]),
    .out(out23)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_115
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[115]),
    .out(out31)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_116
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[116]),
    .out(out39)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_117
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[117]),
    .out(out47)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_118
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[118]),
    .out(out55)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_119
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[119]),
    .out(out63)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_120
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[120]),
    .out(out71)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_121
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[121]),
    .out(out79)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_122
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[122]),
    .out(out87)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_123
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[123]),
    .out(out95)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_124
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[124]),
    .out(out103)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_125
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[125]),
    .out(out111)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_126
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[126]),
    .out(out119)
  );


  reg_pipe
  #(
    .NUM_STAGES(PIPE_EXTRA + 1),
    .DATA_WIDTH(WIDTH)
  )
  reg_in_4_127
  (
    .clk(clk),
    .rst(1'b0),
    .en(en),
    .in(in_reg_wire_7[127]),
    .out(out127)
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_0
  (
    .sel(conf_out[23:0]),
    .in0(in_reg_wire_0[0]),
    .in1(in_reg_wire_0[16]),
    .in2(in_reg_wire_0[32]),
    .in3(in_reg_wire_0[48]),
    .in4(in_reg_wire_0[64]),
    .in5(in_reg_wire_0[80]),
    .in6(in_reg_wire_0[96]),
    .in7(in_reg_wire_0[112]),
    .out0(in_reg_wire_1[0]),
    .out1(in_reg_wire_1[1]),
    .out2(in_reg_wire_1[2]),
    .out3(in_reg_wire_1[3]),
    .out4(in_reg_wire_1[4]),
    .out5(in_reg_wire_1[5]),
    .out6(in_reg_wire_1[6]),
    .out7(in_reg_wire_1[7])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_1
  (
    .sel(conf_out[47:24]),
    .in0(in_reg_wire_0[1]),
    .in1(in_reg_wire_0[17]),
    .in2(in_reg_wire_0[33]),
    .in3(in_reg_wire_0[49]),
    .in4(in_reg_wire_0[65]),
    .in5(in_reg_wire_0[81]),
    .in6(in_reg_wire_0[97]),
    .in7(in_reg_wire_0[113]),
    .out0(in_reg_wire_1[8]),
    .out1(in_reg_wire_1[9]),
    .out2(in_reg_wire_1[10]),
    .out3(in_reg_wire_1[11]),
    .out4(in_reg_wire_1[12]),
    .out5(in_reg_wire_1[13]),
    .out6(in_reg_wire_1[14]),
    .out7(in_reg_wire_1[15])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_2
  (
    .sel(conf_out[71:48]),
    .in0(in_reg_wire_0[2]),
    .in1(in_reg_wire_0[18]),
    .in2(in_reg_wire_0[34]),
    .in3(in_reg_wire_0[50]),
    .in4(in_reg_wire_0[66]),
    .in5(in_reg_wire_0[82]),
    .in6(in_reg_wire_0[98]),
    .in7(in_reg_wire_0[114]),
    .out0(in_reg_wire_1[16]),
    .out1(in_reg_wire_1[17]),
    .out2(in_reg_wire_1[18]),
    .out3(in_reg_wire_1[19]),
    .out4(in_reg_wire_1[20]),
    .out5(in_reg_wire_1[21]),
    .out6(in_reg_wire_1[22]),
    .out7(in_reg_wire_1[23])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_3
  (
    .sel(conf_out[95:72]),
    .in0(in_reg_wire_0[3]),
    .in1(in_reg_wire_0[19]),
    .in2(in_reg_wire_0[35]),
    .in3(in_reg_wire_0[51]),
    .in4(in_reg_wire_0[67]),
    .in5(in_reg_wire_0[83]),
    .in6(in_reg_wire_0[99]),
    .in7(in_reg_wire_0[115]),
    .out0(in_reg_wire_1[24]),
    .out1(in_reg_wire_1[25]),
    .out2(in_reg_wire_1[26]),
    .out3(in_reg_wire_1[27]),
    .out4(in_reg_wire_1[28]),
    .out5(in_reg_wire_1[29]),
    .out6(in_reg_wire_1[30]),
    .out7(in_reg_wire_1[31])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_4
  (
    .sel(conf_out[119:96]),
    .in0(in_reg_wire_0[4]),
    .in1(in_reg_wire_0[20]),
    .in2(in_reg_wire_0[36]),
    .in3(in_reg_wire_0[52]),
    .in4(in_reg_wire_0[68]),
    .in5(in_reg_wire_0[84]),
    .in6(in_reg_wire_0[100]),
    .in7(in_reg_wire_0[116]),
    .out0(in_reg_wire_1[32]),
    .out1(in_reg_wire_1[33]),
    .out2(in_reg_wire_1[34]),
    .out3(in_reg_wire_1[35]),
    .out4(in_reg_wire_1[36]),
    .out5(in_reg_wire_1[37]),
    .out6(in_reg_wire_1[38]),
    .out7(in_reg_wire_1[39])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_5
  (
    .sel(conf_out[143:120]),
    .in0(in_reg_wire_0[5]),
    .in1(in_reg_wire_0[21]),
    .in2(in_reg_wire_0[37]),
    .in3(in_reg_wire_0[53]),
    .in4(in_reg_wire_0[69]),
    .in5(in_reg_wire_0[85]),
    .in6(in_reg_wire_0[101]),
    .in7(in_reg_wire_0[117]),
    .out0(in_reg_wire_1[40]),
    .out1(in_reg_wire_1[41]),
    .out2(in_reg_wire_1[42]),
    .out3(in_reg_wire_1[43]),
    .out4(in_reg_wire_1[44]),
    .out5(in_reg_wire_1[45]),
    .out6(in_reg_wire_1[46]),
    .out7(in_reg_wire_1[47])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_6
  (
    .sel(conf_out[167:144]),
    .in0(in_reg_wire_0[6]),
    .in1(in_reg_wire_0[22]),
    .in2(in_reg_wire_0[38]),
    .in3(in_reg_wire_0[54]),
    .in4(in_reg_wire_0[70]),
    .in5(in_reg_wire_0[86]),
    .in6(in_reg_wire_0[102]),
    .in7(in_reg_wire_0[118]),
    .out0(in_reg_wire_1[48]),
    .out1(in_reg_wire_1[49]),
    .out2(in_reg_wire_1[50]),
    .out3(in_reg_wire_1[51]),
    .out4(in_reg_wire_1[52]),
    .out5(in_reg_wire_1[53]),
    .out6(in_reg_wire_1[54]),
    .out7(in_reg_wire_1[55])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_7
  (
    .sel(conf_out[191:168]),
    .in0(in_reg_wire_0[7]),
    .in1(in_reg_wire_0[23]),
    .in2(in_reg_wire_0[39]),
    .in3(in_reg_wire_0[55]),
    .in4(in_reg_wire_0[71]),
    .in5(in_reg_wire_0[87]),
    .in6(in_reg_wire_0[103]),
    .in7(in_reg_wire_0[119]),
    .out0(in_reg_wire_1[56]),
    .out1(in_reg_wire_1[57]),
    .out2(in_reg_wire_1[58]),
    .out3(in_reg_wire_1[59]),
    .out4(in_reg_wire_1[60]),
    .out5(in_reg_wire_1[61]),
    .out6(in_reg_wire_1[62]),
    .out7(in_reg_wire_1[63])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_8
  (
    .sel(conf_out[215:192]),
    .in0(in_reg_wire_0[8]),
    .in1(in_reg_wire_0[24]),
    .in2(in_reg_wire_0[40]),
    .in3(in_reg_wire_0[56]),
    .in4(in_reg_wire_0[72]),
    .in5(in_reg_wire_0[88]),
    .in6(in_reg_wire_0[104]),
    .in7(in_reg_wire_0[120]),
    .out0(in_reg_wire_1[64]),
    .out1(in_reg_wire_1[65]),
    .out2(in_reg_wire_1[66]),
    .out3(in_reg_wire_1[67]),
    .out4(in_reg_wire_1[68]),
    .out5(in_reg_wire_1[69]),
    .out6(in_reg_wire_1[70]),
    .out7(in_reg_wire_1[71])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_9
  (
    .sel(conf_out[239:216]),
    .in0(in_reg_wire_0[9]),
    .in1(in_reg_wire_0[25]),
    .in2(in_reg_wire_0[41]),
    .in3(in_reg_wire_0[57]),
    .in4(in_reg_wire_0[73]),
    .in5(in_reg_wire_0[89]),
    .in6(in_reg_wire_0[105]),
    .in7(in_reg_wire_0[121]),
    .out0(in_reg_wire_1[72]),
    .out1(in_reg_wire_1[73]),
    .out2(in_reg_wire_1[74]),
    .out3(in_reg_wire_1[75]),
    .out4(in_reg_wire_1[76]),
    .out5(in_reg_wire_1[77]),
    .out6(in_reg_wire_1[78]),
    .out7(in_reg_wire_1[79])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_10
  (
    .sel(conf_out[263:240]),
    .in0(in_reg_wire_0[10]),
    .in1(in_reg_wire_0[26]),
    .in2(in_reg_wire_0[42]),
    .in3(in_reg_wire_0[58]),
    .in4(in_reg_wire_0[74]),
    .in5(in_reg_wire_0[90]),
    .in6(in_reg_wire_0[106]),
    .in7(in_reg_wire_0[122]),
    .out0(in_reg_wire_1[80]),
    .out1(in_reg_wire_1[81]),
    .out2(in_reg_wire_1[82]),
    .out3(in_reg_wire_1[83]),
    .out4(in_reg_wire_1[84]),
    .out5(in_reg_wire_1[85]),
    .out6(in_reg_wire_1[86]),
    .out7(in_reg_wire_1[87])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_11
  (
    .sel(conf_out[287:264]),
    .in0(in_reg_wire_0[11]),
    .in1(in_reg_wire_0[27]),
    .in2(in_reg_wire_0[43]),
    .in3(in_reg_wire_0[59]),
    .in4(in_reg_wire_0[75]),
    .in5(in_reg_wire_0[91]),
    .in6(in_reg_wire_0[107]),
    .in7(in_reg_wire_0[123]),
    .out0(in_reg_wire_1[88]),
    .out1(in_reg_wire_1[89]),
    .out2(in_reg_wire_1[90]),
    .out3(in_reg_wire_1[91]),
    .out4(in_reg_wire_1[92]),
    .out5(in_reg_wire_1[93]),
    .out6(in_reg_wire_1[94]),
    .out7(in_reg_wire_1[95])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_12
  (
    .sel(conf_out[311:288]),
    .in0(in_reg_wire_0[12]),
    .in1(in_reg_wire_0[28]),
    .in2(in_reg_wire_0[44]),
    .in3(in_reg_wire_0[60]),
    .in4(in_reg_wire_0[76]),
    .in5(in_reg_wire_0[92]),
    .in6(in_reg_wire_0[108]),
    .in7(in_reg_wire_0[124]),
    .out0(in_reg_wire_1[96]),
    .out1(in_reg_wire_1[97]),
    .out2(in_reg_wire_1[98]),
    .out3(in_reg_wire_1[99]),
    .out4(in_reg_wire_1[100]),
    .out5(in_reg_wire_1[101]),
    .out6(in_reg_wire_1[102]),
    .out7(in_reg_wire_1[103])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_13
  (
    .sel(conf_out[335:312]),
    .in0(in_reg_wire_0[13]),
    .in1(in_reg_wire_0[29]),
    .in2(in_reg_wire_0[45]),
    .in3(in_reg_wire_0[61]),
    .in4(in_reg_wire_0[77]),
    .in5(in_reg_wire_0[93]),
    .in6(in_reg_wire_0[109]),
    .in7(in_reg_wire_0[125]),
    .out0(in_reg_wire_1[104]),
    .out1(in_reg_wire_1[105]),
    .out2(in_reg_wire_1[106]),
    .out3(in_reg_wire_1[107]),
    .out4(in_reg_wire_1[108]),
    .out5(in_reg_wire_1[109]),
    .out6(in_reg_wire_1[110]),
    .out7(in_reg_wire_1[111])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_14
  (
    .sel(conf_out[359:336]),
    .in0(in_reg_wire_0[14]),
    .in1(in_reg_wire_0[30]),
    .in2(in_reg_wire_0[46]),
    .in3(in_reg_wire_0[62]),
    .in4(in_reg_wire_0[78]),
    .in5(in_reg_wire_0[94]),
    .in6(in_reg_wire_0[110]),
    .in7(in_reg_wire_0[126]),
    .out0(in_reg_wire_1[112]),
    .out1(in_reg_wire_1[113]),
    .out2(in_reg_wire_1[114]),
    .out3(in_reg_wire_1[115]),
    .out4(in_reg_wire_1[116]),
    .out5(in_reg_wire_1[117]),
    .out6(in_reg_wire_1[118]),
    .out7(in_reg_wire_1[119])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_0_15
  (
    .sel(conf_out[383:360]),
    .in0(in_reg_wire_0[15]),
    .in1(in_reg_wire_0[31]),
    .in2(in_reg_wire_0[47]),
    .in3(in_reg_wire_0[63]),
    .in4(in_reg_wire_0[79]),
    .in5(in_reg_wire_0[95]),
    .in6(in_reg_wire_0[111]),
    .in7(in_reg_wire_0[127]),
    .out0(in_reg_wire_1[120]),
    .out1(in_reg_wire_1[121]),
    .out2(in_reg_wire_1[122]),
    .out3(in_reg_wire_1[123]),
    .out4(in_reg_wire_1[124]),
    .out5(in_reg_wire_1[125]),
    .out6(in_reg_wire_1[126]),
    .out7(in_reg_wire_1[127])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_0
  (
    .sel(conf_out[407:384]),
    .in0(in_reg_wire_2[0]),
    .in1(in_reg_wire_2[16]),
    .in2(in_reg_wire_2[32]),
    .in3(in_reg_wire_2[48]),
    .in4(in_reg_wire_2[64]),
    .in5(in_reg_wire_2[80]),
    .in6(in_reg_wire_2[96]),
    .in7(in_reg_wire_2[112]),
    .out0(in_reg_wire_3[0]),
    .out1(in_reg_wire_3[1]),
    .out2(in_reg_wire_3[2]),
    .out3(in_reg_wire_3[3]),
    .out4(in_reg_wire_3[4]),
    .out5(in_reg_wire_3[5]),
    .out6(in_reg_wire_3[6]),
    .out7(in_reg_wire_3[7])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_1
  (
    .sel(conf_out[431:408]),
    .in0(in_reg_wire_2[1]),
    .in1(in_reg_wire_2[17]),
    .in2(in_reg_wire_2[33]),
    .in3(in_reg_wire_2[49]),
    .in4(in_reg_wire_2[65]),
    .in5(in_reg_wire_2[81]),
    .in6(in_reg_wire_2[97]),
    .in7(in_reg_wire_2[113]),
    .out0(in_reg_wire_3[8]),
    .out1(in_reg_wire_3[9]),
    .out2(in_reg_wire_3[10]),
    .out3(in_reg_wire_3[11]),
    .out4(in_reg_wire_3[12]),
    .out5(in_reg_wire_3[13]),
    .out6(in_reg_wire_3[14]),
    .out7(in_reg_wire_3[15])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_2
  (
    .sel(conf_out[455:432]),
    .in0(in_reg_wire_2[2]),
    .in1(in_reg_wire_2[18]),
    .in2(in_reg_wire_2[34]),
    .in3(in_reg_wire_2[50]),
    .in4(in_reg_wire_2[66]),
    .in5(in_reg_wire_2[82]),
    .in6(in_reg_wire_2[98]),
    .in7(in_reg_wire_2[114]),
    .out0(in_reg_wire_3[16]),
    .out1(in_reg_wire_3[17]),
    .out2(in_reg_wire_3[18]),
    .out3(in_reg_wire_3[19]),
    .out4(in_reg_wire_3[20]),
    .out5(in_reg_wire_3[21]),
    .out6(in_reg_wire_3[22]),
    .out7(in_reg_wire_3[23])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_3
  (
    .sel(conf_out[479:456]),
    .in0(in_reg_wire_2[3]),
    .in1(in_reg_wire_2[19]),
    .in2(in_reg_wire_2[35]),
    .in3(in_reg_wire_2[51]),
    .in4(in_reg_wire_2[67]),
    .in5(in_reg_wire_2[83]),
    .in6(in_reg_wire_2[99]),
    .in7(in_reg_wire_2[115]),
    .out0(in_reg_wire_3[24]),
    .out1(in_reg_wire_3[25]),
    .out2(in_reg_wire_3[26]),
    .out3(in_reg_wire_3[27]),
    .out4(in_reg_wire_3[28]),
    .out5(in_reg_wire_3[29]),
    .out6(in_reg_wire_3[30]),
    .out7(in_reg_wire_3[31])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_4
  (
    .sel(conf_out[503:480]),
    .in0(in_reg_wire_2[4]),
    .in1(in_reg_wire_2[20]),
    .in2(in_reg_wire_2[36]),
    .in3(in_reg_wire_2[52]),
    .in4(in_reg_wire_2[68]),
    .in5(in_reg_wire_2[84]),
    .in6(in_reg_wire_2[100]),
    .in7(in_reg_wire_2[116]),
    .out0(in_reg_wire_3[32]),
    .out1(in_reg_wire_3[33]),
    .out2(in_reg_wire_3[34]),
    .out3(in_reg_wire_3[35]),
    .out4(in_reg_wire_3[36]),
    .out5(in_reg_wire_3[37]),
    .out6(in_reg_wire_3[38]),
    .out7(in_reg_wire_3[39])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_5
  (
    .sel(conf_out[527:504]),
    .in0(in_reg_wire_2[5]),
    .in1(in_reg_wire_2[21]),
    .in2(in_reg_wire_2[37]),
    .in3(in_reg_wire_2[53]),
    .in4(in_reg_wire_2[69]),
    .in5(in_reg_wire_2[85]),
    .in6(in_reg_wire_2[101]),
    .in7(in_reg_wire_2[117]),
    .out0(in_reg_wire_3[40]),
    .out1(in_reg_wire_3[41]),
    .out2(in_reg_wire_3[42]),
    .out3(in_reg_wire_3[43]),
    .out4(in_reg_wire_3[44]),
    .out5(in_reg_wire_3[45]),
    .out6(in_reg_wire_3[46]),
    .out7(in_reg_wire_3[47])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_6
  (
    .sel(conf_out[551:528]),
    .in0(in_reg_wire_2[6]),
    .in1(in_reg_wire_2[22]),
    .in2(in_reg_wire_2[38]),
    .in3(in_reg_wire_2[54]),
    .in4(in_reg_wire_2[70]),
    .in5(in_reg_wire_2[86]),
    .in6(in_reg_wire_2[102]),
    .in7(in_reg_wire_2[118]),
    .out0(in_reg_wire_3[48]),
    .out1(in_reg_wire_3[49]),
    .out2(in_reg_wire_3[50]),
    .out3(in_reg_wire_3[51]),
    .out4(in_reg_wire_3[52]),
    .out5(in_reg_wire_3[53]),
    .out6(in_reg_wire_3[54]),
    .out7(in_reg_wire_3[55])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_7
  (
    .sel(conf_out[575:552]),
    .in0(in_reg_wire_2[7]),
    .in1(in_reg_wire_2[23]),
    .in2(in_reg_wire_2[39]),
    .in3(in_reg_wire_2[55]),
    .in4(in_reg_wire_2[71]),
    .in5(in_reg_wire_2[87]),
    .in6(in_reg_wire_2[103]),
    .in7(in_reg_wire_2[119]),
    .out0(in_reg_wire_3[56]),
    .out1(in_reg_wire_3[57]),
    .out2(in_reg_wire_3[58]),
    .out3(in_reg_wire_3[59]),
    .out4(in_reg_wire_3[60]),
    .out5(in_reg_wire_3[61]),
    .out6(in_reg_wire_3[62]),
    .out7(in_reg_wire_3[63])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_8
  (
    .sel(conf_out[599:576]),
    .in0(in_reg_wire_2[8]),
    .in1(in_reg_wire_2[24]),
    .in2(in_reg_wire_2[40]),
    .in3(in_reg_wire_2[56]),
    .in4(in_reg_wire_2[72]),
    .in5(in_reg_wire_2[88]),
    .in6(in_reg_wire_2[104]),
    .in7(in_reg_wire_2[120]),
    .out0(in_reg_wire_3[64]),
    .out1(in_reg_wire_3[65]),
    .out2(in_reg_wire_3[66]),
    .out3(in_reg_wire_3[67]),
    .out4(in_reg_wire_3[68]),
    .out5(in_reg_wire_3[69]),
    .out6(in_reg_wire_3[70]),
    .out7(in_reg_wire_3[71])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_9
  (
    .sel(conf_out[623:600]),
    .in0(in_reg_wire_2[9]),
    .in1(in_reg_wire_2[25]),
    .in2(in_reg_wire_2[41]),
    .in3(in_reg_wire_2[57]),
    .in4(in_reg_wire_2[73]),
    .in5(in_reg_wire_2[89]),
    .in6(in_reg_wire_2[105]),
    .in7(in_reg_wire_2[121]),
    .out0(in_reg_wire_3[72]),
    .out1(in_reg_wire_3[73]),
    .out2(in_reg_wire_3[74]),
    .out3(in_reg_wire_3[75]),
    .out4(in_reg_wire_3[76]),
    .out5(in_reg_wire_3[77]),
    .out6(in_reg_wire_3[78]),
    .out7(in_reg_wire_3[79])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_10
  (
    .sel(conf_out[647:624]),
    .in0(in_reg_wire_2[10]),
    .in1(in_reg_wire_2[26]),
    .in2(in_reg_wire_2[42]),
    .in3(in_reg_wire_2[58]),
    .in4(in_reg_wire_2[74]),
    .in5(in_reg_wire_2[90]),
    .in6(in_reg_wire_2[106]),
    .in7(in_reg_wire_2[122]),
    .out0(in_reg_wire_3[80]),
    .out1(in_reg_wire_3[81]),
    .out2(in_reg_wire_3[82]),
    .out3(in_reg_wire_3[83]),
    .out4(in_reg_wire_3[84]),
    .out5(in_reg_wire_3[85]),
    .out6(in_reg_wire_3[86]),
    .out7(in_reg_wire_3[87])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_11
  (
    .sel(conf_out[671:648]),
    .in0(in_reg_wire_2[11]),
    .in1(in_reg_wire_2[27]),
    .in2(in_reg_wire_2[43]),
    .in3(in_reg_wire_2[59]),
    .in4(in_reg_wire_2[75]),
    .in5(in_reg_wire_2[91]),
    .in6(in_reg_wire_2[107]),
    .in7(in_reg_wire_2[123]),
    .out0(in_reg_wire_3[88]),
    .out1(in_reg_wire_3[89]),
    .out2(in_reg_wire_3[90]),
    .out3(in_reg_wire_3[91]),
    .out4(in_reg_wire_3[92]),
    .out5(in_reg_wire_3[93]),
    .out6(in_reg_wire_3[94]),
    .out7(in_reg_wire_3[95])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_12
  (
    .sel(conf_out[695:672]),
    .in0(in_reg_wire_2[12]),
    .in1(in_reg_wire_2[28]),
    .in2(in_reg_wire_2[44]),
    .in3(in_reg_wire_2[60]),
    .in4(in_reg_wire_2[76]),
    .in5(in_reg_wire_2[92]),
    .in6(in_reg_wire_2[108]),
    .in7(in_reg_wire_2[124]),
    .out0(in_reg_wire_3[96]),
    .out1(in_reg_wire_3[97]),
    .out2(in_reg_wire_3[98]),
    .out3(in_reg_wire_3[99]),
    .out4(in_reg_wire_3[100]),
    .out5(in_reg_wire_3[101]),
    .out6(in_reg_wire_3[102]),
    .out7(in_reg_wire_3[103])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_13
  (
    .sel(conf_out[719:696]),
    .in0(in_reg_wire_2[13]),
    .in1(in_reg_wire_2[29]),
    .in2(in_reg_wire_2[45]),
    .in3(in_reg_wire_2[61]),
    .in4(in_reg_wire_2[77]),
    .in5(in_reg_wire_2[93]),
    .in6(in_reg_wire_2[109]),
    .in7(in_reg_wire_2[125]),
    .out0(in_reg_wire_3[104]),
    .out1(in_reg_wire_3[105]),
    .out2(in_reg_wire_3[106]),
    .out3(in_reg_wire_3[107]),
    .out4(in_reg_wire_3[108]),
    .out5(in_reg_wire_3[109]),
    .out6(in_reg_wire_3[110]),
    .out7(in_reg_wire_3[111])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_14
  (
    .sel(conf_out[743:720]),
    .in0(in_reg_wire_2[14]),
    .in1(in_reg_wire_2[30]),
    .in2(in_reg_wire_2[46]),
    .in3(in_reg_wire_2[62]),
    .in4(in_reg_wire_2[78]),
    .in5(in_reg_wire_2[94]),
    .in6(in_reg_wire_2[110]),
    .in7(in_reg_wire_2[126]),
    .out0(in_reg_wire_3[112]),
    .out1(in_reg_wire_3[113]),
    .out2(in_reg_wire_3[114]),
    .out3(in_reg_wire_3[115]),
    .out4(in_reg_wire_3[116]),
    .out5(in_reg_wire_3[117]),
    .out6(in_reg_wire_3[118]),
    .out7(in_reg_wire_3[119])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_1_15
  (
    .sel(conf_out[767:744]),
    .in0(in_reg_wire_2[15]),
    .in1(in_reg_wire_2[31]),
    .in2(in_reg_wire_2[47]),
    .in3(in_reg_wire_2[63]),
    .in4(in_reg_wire_2[79]),
    .in5(in_reg_wire_2[95]),
    .in6(in_reg_wire_2[111]),
    .in7(in_reg_wire_2[127]),
    .out0(in_reg_wire_3[120]),
    .out1(in_reg_wire_3[121]),
    .out2(in_reg_wire_3[122]),
    .out3(in_reg_wire_3[123]),
    .out4(in_reg_wire_3[124]),
    .out5(in_reg_wire_3[125]),
    .out6(in_reg_wire_3[126]),
    .out7(in_reg_wire_3[127])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_0
  (
    .sel(conf_out[791:768]),
    .in0(in_reg_wire_4[0]),
    .in1(in_reg_wire_4[16]),
    .in2(in_reg_wire_4[32]),
    .in3(in_reg_wire_4[48]),
    .in4(in_reg_wire_4[64]),
    .in5(in_reg_wire_4[80]),
    .in6(in_reg_wire_4[96]),
    .in7(in_reg_wire_4[112]),
    .out0(in_reg_wire_5[0]),
    .out1(in_reg_wire_5[1]),
    .out2(in_reg_wire_5[2]),
    .out3(in_reg_wire_5[3]),
    .out4(in_reg_wire_5[4]),
    .out5(in_reg_wire_5[5]),
    .out6(in_reg_wire_5[6]),
    .out7(in_reg_wire_5[7])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_1
  (
    .sel(conf_out[815:792]),
    .in0(in_reg_wire_4[1]),
    .in1(in_reg_wire_4[17]),
    .in2(in_reg_wire_4[33]),
    .in3(in_reg_wire_4[49]),
    .in4(in_reg_wire_4[65]),
    .in5(in_reg_wire_4[81]),
    .in6(in_reg_wire_4[97]),
    .in7(in_reg_wire_4[113]),
    .out0(in_reg_wire_5[8]),
    .out1(in_reg_wire_5[9]),
    .out2(in_reg_wire_5[10]),
    .out3(in_reg_wire_5[11]),
    .out4(in_reg_wire_5[12]),
    .out5(in_reg_wire_5[13]),
    .out6(in_reg_wire_5[14]),
    .out7(in_reg_wire_5[15])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_2
  (
    .sel(conf_out[839:816]),
    .in0(in_reg_wire_4[2]),
    .in1(in_reg_wire_4[18]),
    .in2(in_reg_wire_4[34]),
    .in3(in_reg_wire_4[50]),
    .in4(in_reg_wire_4[66]),
    .in5(in_reg_wire_4[82]),
    .in6(in_reg_wire_4[98]),
    .in7(in_reg_wire_4[114]),
    .out0(in_reg_wire_5[16]),
    .out1(in_reg_wire_5[17]),
    .out2(in_reg_wire_5[18]),
    .out3(in_reg_wire_5[19]),
    .out4(in_reg_wire_5[20]),
    .out5(in_reg_wire_5[21]),
    .out6(in_reg_wire_5[22]),
    .out7(in_reg_wire_5[23])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_3
  (
    .sel(conf_out[863:840]),
    .in0(in_reg_wire_4[3]),
    .in1(in_reg_wire_4[19]),
    .in2(in_reg_wire_4[35]),
    .in3(in_reg_wire_4[51]),
    .in4(in_reg_wire_4[67]),
    .in5(in_reg_wire_4[83]),
    .in6(in_reg_wire_4[99]),
    .in7(in_reg_wire_4[115]),
    .out0(in_reg_wire_5[24]),
    .out1(in_reg_wire_5[25]),
    .out2(in_reg_wire_5[26]),
    .out3(in_reg_wire_5[27]),
    .out4(in_reg_wire_5[28]),
    .out5(in_reg_wire_5[29]),
    .out6(in_reg_wire_5[30]),
    .out7(in_reg_wire_5[31])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_4
  (
    .sel(conf_out[887:864]),
    .in0(in_reg_wire_4[4]),
    .in1(in_reg_wire_4[20]),
    .in2(in_reg_wire_4[36]),
    .in3(in_reg_wire_4[52]),
    .in4(in_reg_wire_4[68]),
    .in5(in_reg_wire_4[84]),
    .in6(in_reg_wire_4[100]),
    .in7(in_reg_wire_4[116]),
    .out0(in_reg_wire_5[32]),
    .out1(in_reg_wire_5[33]),
    .out2(in_reg_wire_5[34]),
    .out3(in_reg_wire_5[35]),
    .out4(in_reg_wire_5[36]),
    .out5(in_reg_wire_5[37]),
    .out6(in_reg_wire_5[38]),
    .out7(in_reg_wire_5[39])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_5
  (
    .sel(conf_out[911:888]),
    .in0(in_reg_wire_4[5]),
    .in1(in_reg_wire_4[21]),
    .in2(in_reg_wire_4[37]),
    .in3(in_reg_wire_4[53]),
    .in4(in_reg_wire_4[69]),
    .in5(in_reg_wire_4[85]),
    .in6(in_reg_wire_4[101]),
    .in7(in_reg_wire_4[117]),
    .out0(in_reg_wire_5[40]),
    .out1(in_reg_wire_5[41]),
    .out2(in_reg_wire_5[42]),
    .out3(in_reg_wire_5[43]),
    .out4(in_reg_wire_5[44]),
    .out5(in_reg_wire_5[45]),
    .out6(in_reg_wire_5[46]),
    .out7(in_reg_wire_5[47])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_6
  (
    .sel(conf_out[935:912]),
    .in0(in_reg_wire_4[6]),
    .in1(in_reg_wire_4[22]),
    .in2(in_reg_wire_4[38]),
    .in3(in_reg_wire_4[54]),
    .in4(in_reg_wire_4[70]),
    .in5(in_reg_wire_4[86]),
    .in6(in_reg_wire_4[102]),
    .in7(in_reg_wire_4[118]),
    .out0(in_reg_wire_5[48]),
    .out1(in_reg_wire_5[49]),
    .out2(in_reg_wire_5[50]),
    .out3(in_reg_wire_5[51]),
    .out4(in_reg_wire_5[52]),
    .out5(in_reg_wire_5[53]),
    .out6(in_reg_wire_5[54]),
    .out7(in_reg_wire_5[55])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_7
  (
    .sel(conf_out[959:936]),
    .in0(in_reg_wire_4[7]),
    .in1(in_reg_wire_4[23]),
    .in2(in_reg_wire_4[39]),
    .in3(in_reg_wire_4[55]),
    .in4(in_reg_wire_4[71]),
    .in5(in_reg_wire_4[87]),
    .in6(in_reg_wire_4[103]),
    .in7(in_reg_wire_4[119]),
    .out0(in_reg_wire_5[56]),
    .out1(in_reg_wire_5[57]),
    .out2(in_reg_wire_5[58]),
    .out3(in_reg_wire_5[59]),
    .out4(in_reg_wire_5[60]),
    .out5(in_reg_wire_5[61]),
    .out6(in_reg_wire_5[62]),
    .out7(in_reg_wire_5[63])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_8
  (
    .sel(conf_out[983:960]),
    .in0(in_reg_wire_4[8]),
    .in1(in_reg_wire_4[24]),
    .in2(in_reg_wire_4[40]),
    .in3(in_reg_wire_4[56]),
    .in4(in_reg_wire_4[72]),
    .in5(in_reg_wire_4[88]),
    .in6(in_reg_wire_4[104]),
    .in7(in_reg_wire_4[120]),
    .out0(in_reg_wire_5[64]),
    .out1(in_reg_wire_5[65]),
    .out2(in_reg_wire_5[66]),
    .out3(in_reg_wire_5[67]),
    .out4(in_reg_wire_5[68]),
    .out5(in_reg_wire_5[69]),
    .out6(in_reg_wire_5[70]),
    .out7(in_reg_wire_5[71])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_9
  (
    .sel(conf_out[1007:984]),
    .in0(in_reg_wire_4[9]),
    .in1(in_reg_wire_4[25]),
    .in2(in_reg_wire_4[41]),
    .in3(in_reg_wire_4[57]),
    .in4(in_reg_wire_4[73]),
    .in5(in_reg_wire_4[89]),
    .in6(in_reg_wire_4[105]),
    .in7(in_reg_wire_4[121]),
    .out0(in_reg_wire_5[72]),
    .out1(in_reg_wire_5[73]),
    .out2(in_reg_wire_5[74]),
    .out3(in_reg_wire_5[75]),
    .out4(in_reg_wire_5[76]),
    .out5(in_reg_wire_5[77]),
    .out6(in_reg_wire_5[78]),
    .out7(in_reg_wire_5[79])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_10
  (
    .sel(conf_out[1031:1008]),
    .in0(in_reg_wire_4[10]),
    .in1(in_reg_wire_4[26]),
    .in2(in_reg_wire_4[42]),
    .in3(in_reg_wire_4[58]),
    .in4(in_reg_wire_4[74]),
    .in5(in_reg_wire_4[90]),
    .in6(in_reg_wire_4[106]),
    .in7(in_reg_wire_4[122]),
    .out0(in_reg_wire_5[80]),
    .out1(in_reg_wire_5[81]),
    .out2(in_reg_wire_5[82]),
    .out3(in_reg_wire_5[83]),
    .out4(in_reg_wire_5[84]),
    .out5(in_reg_wire_5[85]),
    .out6(in_reg_wire_5[86]),
    .out7(in_reg_wire_5[87])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_11
  (
    .sel(conf_out[1055:1032]),
    .in0(in_reg_wire_4[11]),
    .in1(in_reg_wire_4[27]),
    .in2(in_reg_wire_4[43]),
    .in3(in_reg_wire_4[59]),
    .in4(in_reg_wire_4[75]),
    .in5(in_reg_wire_4[91]),
    .in6(in_reg_wire_4[107]),
    .in7(in_reg_wire_4[123]),
    .out0(in_reg_wire_5[88]),
    .out1(in_reg_wire_5[89]),
    .out2(in_reg_wire_5[90]),
    .out3(in_reg_wire_5[91]),
    .out4(in_reg_wire_5[92]),
    .out5(in_reg_wire_5[93]),
    .out6(in_reg_wire_5[94]),
    .out7(in_reg_wire_5[95])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_12
  (
    .sel(conf_out[1079:1056]),
    .in0(in_reg_wire_4[12]),
    .in1(in_reg_wire_4[28]),
    .in2(in_reg_wire_4[44]),
    .in3(in_reg_wire_4[60]),
    .in4(in_reg_wire_4[76]),
    .in5(in_reg_wire_4[92]),
    .in6(in_reg_wire_4[108]),
    .in7(in_reg_wire_4[124]),
    .out0(in_reg_wire_5[96]),
    .out1(in_reg_wire_5[97]),
    .out2(in_reg_wire_5[98]),
    .out3(in_reg_wire_5[99]),
    .out4(in_reg_wire_5[100]),
    .out5(in_reg_wire_5[101]),
    .out6(in_reg_wire_5[102]),
    .out7(in_reg_wire_5[103])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_13
  (
    .sel(conf_out[1103:1080]),
    .in0(in_reg_wire_4[13]),
    .in1(in_reg_wire_4[29]),
    .in2(in_reg_wire_4[45]),
    .in3(in_reg_wire_4[61]),
    .in4(in_reg_wire_4[77]),
    .in5(in_reg_wire_4[93]),
    .in6(in_reg_wire_4[109]),
    .in7(in_reg_wire_4[125]),
    .out0(in_reg_wire_5[104]),
    .out1(in_reg_wire_5[105]),
    .out2(in_reg_wire_5[106]),
    .out3(in_reg_wire_5[107]),
    .out4(in_reg_wire_5[108]),
    .out5(in_reg_wire_5[109]),
    .out6(in_reg_wire_5[110]),
    .out7(in_reg_wire_5[111])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_14
  (
    .sel(conf_out[1127:1104]),
    .in0(in_reg_wire_4[14]),
    .in1(in_reg_wire_4[30]),
    .in2(in_reg_wire_4[46]),
    .in3(in_reg_wire_4[62]),
    .in4(in_reg_wire_4[78]),
    .in5(in_reg_wire_4[94]),
    .in6(in_reg_wire_4[110]),
    .in7(in_reg_wire_4[126]),
    .out0(in_reg_wire_5[112]),
    .out1(in_reg_wire_5[113]),
    .out2(in_reg_wire_5[114]),
    .out3(in_reg_wire_5[115]),
    .out4(in_reg_wire_5[116]),
    .out5(in_reg_wire_5[117]),
    .out6(in_reg_wire_5[118]),
    .out7(in_reg_wire_5[119])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_2_15
  (
    .sel(conf_out[1151:1128]),
    .in0(in_reg_wire_4[15]),
    .in1(in_reg_wire_4[31]),
    .in2(in_reg_wire_4[47]),
    .in3(in_reg_wire_4[63]),
    .in4(in_reg_wire_4[79]),
    .in5(in_reg_wire_4[95]),
    .in6(in_reg_wire_4[111]),
    .in7(in_reg_wire_4[127]),
    .out0(in_reg_wire_5[120]),
    .out1(in_reg_wire_5[121]),
    .out2(in_reg_wire_5[122]),
    .out3(in_reg_wire_5[123]),
    .out4(in_reg_wire_5[124]),
    .out5(in_reg_wire_5[125]),
    .out6(in_reg_wire_5[126]),
    .out7(in_reg_wire_5[127])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_3_0
  (
    .sel(conf_out[1175:1152]),
    .in0(in_reg_wire_6[0]),
    .in1(in_reg_wire_6[16]),
    .in2(in_reg_wire_6[32]),
    .in3(in_reg_wire_6[48]),
    .in4(in_reg_wire_6[64]),
    .in5(in_reg_wire_6[80]),
    .in6(in_reg_wire_6[96]),
    .in7(in_reg_wire_6[112]),
    .out0(in_reg_wire_7[0]),
    .out1(in_reg_wire_7[1]),
    .out2(in_reg_wire_7[2]),
    .out3(in_reg_wire_7[3]),
    .out4(in_reg_wire_7[4]),
    .out5(in_reg_wire_7[5]),
    .out6(in_reg_wire_7[6]),
    .out7(in_reg_wire_7[7])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_3_1
  (
    .sel(conf_out[1199:1176]),
    .in0(in_reg_wire_6[1]),
    .in1(in_reg_wire_6[17]),
    .in2(in_reg_wire_6[33]),
    .in3(in_reg_wire_6[49]),
    .in4(in_reg_wire_6[65]),
    .in5(in_reg_wire_6[81]),
    .in6(in_reg_wire_6[97]),
    .in7(in_reg_wire_6[113]),
    .out0(in_reg_wire_7[8]),
    .out1(in_reg_wire_7[9]),
    .out2(in_reg_wire_7[10]),
    .out3(in_reg_wire_7[11]),
    .out4(in_reg_wire_7[12]),
    .out5(in_reg_wire_7[13]),
    .out6(in_reg_wire_7[14]),
    .out7(in_reg_wire_7[15])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_3_2
  (
    .sel(conf_out[1223:1200]),
    .in0(in_reg_wire_6[2]),
    .in1(in_reg_wire_6[18]),
    .in2(in_reg_wire_6[34]),
    .in3(in_reg_wire_6[50]),
    .in4(in_reg_wire_6[66]),
    .in5(in_reg_wire_6[82]),
    .in6(in_reg_wire_6[98]),
    .in7(in_reg_wire_6[114]),
    .out0(in_reg_wire_7[16]),
    .out1(in_reg_wire_7[17]),
    .out2(in_reg_wire_7[18]),
    .out3(in_reg_wire_7[19]),
    .out4(in_reg_wire_7[20]),
    .out5(in_reg_wire_7[21]),
    .out6(in_reg_wire_7[22]),
    .out7(in_reg_wire_7[23])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_3_3
  (
    .sel(conf_out[1247:1224]),
    .in0(in_reg_wire_6[3]),
    .in1(in_reg_wire_6[19]),
    .in2(in_reg_wire_6[35]),
    .in3(in_reg_wire_6[51]),
    .in4(in_reg_wire_6[67]),
    .in5(in_reg_wire_6[83]),
    .in6(in_reg_wire_6[99]),
    .in7(in_reg_wire_6[115]),
    .out0(in_reg_wire_7[24]),
    .out1(in_reg_wire_7[25]),
    .out2(in_reg_wire_7[26]),
    .out3(in_reg_wire_7[27]),
    .out4(in_reg_wire_7[28]),
    .out5(in_reg_wire_7[29]),
    .out6(in_reg_wire_7[30]),
    .out7(in_reg_wire_7[31])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_3_4
  (
    .sel(conf_out[1271:1248]),
    .in0(in_reg_wire_6[4]),
    .in1(in_reg_wire_6[20]),
    .in2(in_reg_wire_6[36]),
    .in3(in_reg_wire_6[52]),
    .in4(in_reg_wire_6[68]),
    .in5(in_reg_wire_6[84]),
    .in6(in_reg_wire_6[100]),
    .in7(in_reg_wire_6[116]),
    .out0(in_reg_wire_7[32]),
    .out1(in_reg_wire_7[33]),
    .out2(in_reg_wire_7[34]),
    .out3(in_reg_wire_7[35]),
    .out4(in_reg_wire_7[36]),
    .out5(in_reg_wire_7[37]),
    .out6(in_reg_wire_7[38]),
    .out7(in_reg_wire_7[39])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_3_5
  (
    .sel(conf_out[1295:1272]),
    .in0(in_reg_wire_6[5]),
    .in1(in_reg_wire_6[21]),
    .in2(in_reg_wire_6[37]),
    .in3(in_reg_wire_6[53]),
    .in4(in_reg_wire_6[69]),
    .in5(in_reg_wire_6[85]),
    .in6(in_reg_wire_6[101]),
    .in7(in_reg_wire_6[117]),
    .out0(in_reg_wire_7[40]),
    .out1(in_reg_wire_7[41]),
    .out2(in_reg_wire_7[42]),
    .out3(in_reg_wire_7[43]),
    .out4(in_reg_wire_7[44]),
    .out5(in_reg_wire_7[45]),
    .out6(in_reg_wire_7[46]),
    .out7(in_reg_wire_7[47])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_3_6
  (
    .sel(conf_out[1319:1296]),
    .in0(in_reg_wire_6[6]),
    .in1(in_reg_wire_6[22]),
    .in2(in_reg_wire_6[38]),
    .in3(in_reg_wire_6[54]),
    .in4(in_reg_wire_6[70]),
    .in5(in_reg_wire_6[86]),
    .in6(in_reg_wire_6[102]),
    .in7(in_reg_wire_6[118]),
    .out0(in_reg_wire_7[48]),
    .out1(in_reg_wire_7[49]),
    .out2(in_reg_wire_7[50]),
    .out3(in_reg_wire_7[51]),
    .out4(in_reg_wire_7[52]),
    .out5(in_reg_wire_7[53]),
    .out6(in_reg_wire_7[54]),
    .out7(in_reg_wire_7[55])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_3_7
  (
    .sel(conf_out[1343:1320]),
    .in0(in_reg_wire_6[7]),
    .in1(in_reg_wire_6[23]),
    .in2(in_reg_wire_6[39]),
    .in3(in_reg_wire_6[55]),
    .in4(in_reg_wire_6[71]),
    .in5(in_reg_wire_6[87]),
    .in6(in_reg_wire_6[103]),
    .in7(in_reg_wire_6[119]),
    .out0(in_reg_wire_7[56]),
    .out1(in_reg_wire_7[57]),
    .out2(in_reg_wire_7[58]),
    .out3(in_reg_wire_7[59]),
    .out4(in_reg_wire_7[60]),
    .out5(in_reg_wire_7[61]),
    .out6(in_reg_wire_7[62]),
    .out7(in_reg_wire_7[63])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_3_8
  (
    .sel(conf_out[1367:1344]),
    .in0(in_reg_wire_6[8]),
    .in1(in_reg_wire_6[24]),
    .in2(in_reg_wire_6[40]),
    .in3(in_reg_wire_6[56]),
    .in4(in_reg_wire_6[72]),
    .in5(in_reg_wire_6[88]),
    .in6(in_reg_wire_6[104]),
    .in7(in_reg_wire_6[120]),
    .out0(in_reg_wire_7[64]),
    .out1(in_reg_wire_7[65]),
    .out2(in_reg_wire_7[66]),
    .out3(in_reg_wire_7[67]),
    .out4(in_reg_wire_7[68]),
    .out5(in_reg_wire_7[69]),
    .out6(in_reg_wire_7[70]),
    .out7(in_reg_wire_7[71])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_3_9
  (
    .sel(conf_out[1391:1368]),
    .in0(in_reg_wire_6[9]),
    .in1(in_reg_wire_6[25]),
    .in2(in_reg_wire_6[41]),
    .in3(in_reg_wire_6[57]),
    .in4(in_reg_wire_6[73]),
    .in5(in_reg_wire_6[89]),
    .in6(in_reg_wire_6[105]),
    .in7(in_reg_wire_6[121]),
    .out0(in_reg_wire_7[72]),
    .out1(in_reg_wire_7[73]),
    .out2(in_reg_wire_7[74]),
    .out3(in_reg_wire_7[75]),
    .out4(in_reg_wire_7[76]),
    .out5(in_reg_wire_7[77]),
    .out6(in_reg_wire_7[78]),
    .out7(in_reg_wire_7[79])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_3_10
  (
    .sel(conf_out[1415:1392]),
    .in0(in_reg_wire_6[10]),
    .in1(in_reg_wire_6[26]),
    .in2(in_reg_wire_6[42]),
    .in3(in_reg_wire_6[58]),
    .in4(in_reg_wire_6[74]),
    .in5(in_reg_wire_6[90]),
    .in6(in_reg_wire_6[106]),
    .in7(in_reg_wire_6[122]),
    .out0(in_reg_wire_7[80]),
    .out1(in_reg_wire_7[81]),
    .out2(in_reg_wire_7[82]),
    .out3(in_reg_wire_7[83]),
    .out4(in_reg_wire_7[84]),
    .out5(in_reg_wire_7[85]),
    .out6(in_reg_wire_7[86]),
    .out7(in_reg_wire_7[87])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_3_11
  (
    .sel(conf_out[1439:1416]),
    .in0(in_reg_wire_6[11]),
    .in1(in_reg_wire_6[27]),
    .in2(in_reg_wire_6[43]),
    .in3(in_reg_wire_6[59]),
    .in4(in_reg_wire_6[75]),
    .in5(in_reg_wire_6[91]),
    .in6(in_reg_wire_6[107]),
    .in7(in_reg_wire_6[123]),
    .out0(in_reg_wire_7[88]),
    .out1(in_reg_wire_7[89]),
    .out2(in_reg_wire_7[90]),
    .out3(in_reg_wire_7[91]),
    .out4(in_reg_wire_7[92]),
    .out5(in_reg_wire_7[93]),
    .out6(in_reg_wire_7[94]),
    .out7(in_reg_wire_7[95])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_3_12
  (
    .sel(conf_out[1463:1440]),
    .in0(in_reg_wire_6[12]),
    .in1(in_reg_wire_6[28]),
    .in2(in_reg_wire_6[44]),
    .in3(in_reg_wire_6[60]),
    .in4(in_reg_wire_6[76]),
    .in5(in_reg_wire_6[92]),
    .in6(in_reg_wire_6[108]),
    .in7(in_reg_wire_6[124]),
    .out0(in_reg_wire_7[96]),
    .out1(in_reg_wire_7[97]),
    .out2(in_reg_wire_7[98]),
    .out3(in_reg_wire_7[99]),
    .out4(in_reg_wire_7[100]),
    .out5(in_reg_wire_7[101]),
    .out6(in_reg_wire_7[102]),
    .out7(in_reg_wire_7[103])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_3_13
  (
    .sel(conf_out[1487:1464]),
    .in0(in_reg_wire_6[13]),
    .in1(in_reg_wire_6[29]),
    .in2(in_reg_wire_6[45]),
    .in3(in_reg_wire_6[61]),
    .in4(in_reg_wire_6[77]),
    .in5(in_reg_wire_6[93]),
    .in6(in_reg_wire_6[109]),
    .in7(in_reg_wire_6[125]),
    .out0(in_reg_wire_7[104]),
    .out1(in_reg_wire_7[105]),
    .out2(in_reg_wire_7[106]),
    .out3(in_reg_wire_7[107]),
    .out4(in_reg_wire_7[108]),
    .out5(in_reg_wire_7[109]),
    .out6(in_reg_wire_7[110]),
    .out7(in_reg_wire_7[111])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_3_14
  (
    .sel(conf_out[1511:1488]),
    .in0(in_reg_wire_6[14]),
    .in1(in_reg_wire_6[30]),
    .in2(in_reg_wire_6[46]),
    .in3(in_reg_wire_6[62]),
    .in4(in_reg_wire_6[78]),
    .in5(in_reg_wire_6[94]),
    .in6(in_reg_wire_6[110]),
    .in7(in_reg_wire_6[126]),
    .out0(in_reg_wire_7[112]),
    .out1(in_reg_wire_7[113]),
    .out2(in_reg_wire_7[114]),
    .out3(in_reg_wire_7[115]),
    .out4(in_reg_wire_7[116]),
    .out5(in_reg_wire_7[117]),
    .out6(in_reg_wire_7[118]),
    .out7(in_reg_wire_7[119])
  );


  switch_box8x8
  #(
    .WIDTH(WIDTH)
  )
  sw_3_15
  (
    .sel(conf_out[1535:1512]),
    .in0(in_reg_wire_6[15]),
    .in1(in_reg_wire_6[31]),
    .in2(in_reg_wire_6[47]),
    .in3(in_reg_wire_6[63]),
    .in4(in_reg_wire_6[79]),
    .in5(in_reg_wire_6[95]),
    .in6(in_reg_wire_6[111]),
    .in7(in_reg_wire_6[127]),
    .out0(in_reg_wire_7[120]),
    .out1(in_reg_wire_7[121]),
    .out2(in_reg_wire_7[122]),
    .out3(in_reg_wire_7[123]),
    .out4(in_reg_wire_7[124]),
    .out5(in_reg_wire_7[125]),
    .out6(in_reg_wire_7[126]),
    .out7(in_reg_wire_7[127])
  );

endmodule